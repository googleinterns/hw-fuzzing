module DUT(
  input         clock,
  input         reset,
  input         io_meta_reset,
  input  [34:0] io_inputs,
  output        io_coverage_0,
  output        io_coverage_1,
  output        io_coverage_2,
  output        io_coverage_3,
  output        io_coverage_4,
  output        io_coverage_5,
  output        io_coverage_6,
  output        io_coverage_7,
  output        io_coverage_8,
  output        io_coverage_9,
  output        io_coverage_10,
  output        io_coverage_11,
  output        io_coverage_12,
  output        io_coverage_13,
  output        io_coverage_14,
  output        io_coverage_15,
  output        io_coverage_16,
  output        io_coverage_17,
  output        io_coverage_18,
  output        io_coverage_19,
  output        io_coverage_20,
  output        io_coverage_21,
  output        io_coverage_22,
  output        io_coverage_23,
  output        io_coverage_24,
  output        io_coverage_25,
  output        io_coverage_26,
  output        io_coverage_27,
  output        io_coverage_28,
  output        io_coverage_29,
  output        io_coverage_30,
  output        io_coverage_31,
  output        io_coverage_32,
  output        io_coverage_33,
  output        io_coverage_34,
  output        io_coverage_35,
  output        io_coverage_36,
  output        io_coverage_37,
  output        io_coverage_38,
  output        io_coverage_39,
  output        io_coverage_40,
  output        io_coverage_41,
  output        io_coverage_42,
  output        io_coverage_43,
  output        io_coverage_44,
  output        io_coverage_45,
  output        io_coverage_46,
  output        io_coverage_47,
  output        io_coverage_48,
  output        io_coverage_49,
  output        io_coverage_50,
  output        io_coverage_51,
  output        io_coverage_52,
  output        io_coverage_53,
  output        io_coverage_54,
  output        io_coverage_55,
  output        io_coverage_56,
  output        io_coverage_57,
  output        io_coverage_58,
  output        io_coverage_59,
  output        io_coverage_60,
  output        io_coverage_61,
  output        io_coverage_62,
  output        io_coverage_63,
  output        io_coverage_64,
  output        io_coverage_65,
  output        io_coverage_66,
  output        io_coverage_67,
  output        io_coverage_68,
  output        io_coverage_69,
  output        io_coverage_70,
  output        io_coverage_71,
  output        io_coverage_72,
  output        io_coverage_73,
  output        io_coverage_74,
  output        io_coverage_75,
  output        io_coverage_76,
  output        io_coverage_77,
  output        io_coverage_78,
  output        io_coverage_79,
  output        io_coverage_80,
  output        io_coverage_81,
  output        io_coverage_82,
  output        io_coverage_83,
  output        io_coverage_84,
  output        io_coverage_85,
  output        io_coverage_86,
  output        io_coverage_87,
  output        io_coverage_88,
  output        io_coverage_89,
  output        io_coverage_90,
  output        io_coverage_91,
  output        io_coverage_92,
  output        io_coverage_93,
  output        io_coverage_94,
  output        io_coverage_95,
  output        io_coverage_96,
  output        io_coverage_97,
  output        io_coverage_98,
  output        io_coverage_99,
  output        io_coverage_100,
  output        io_coverage_101,
  output        io_coverage_102,
  output        io_coverage_103,
  output        io_coverage_104,
  output        io_coverage_105,
  output        io_coverage_106,
  output        io_coverage_107,
  output        io_coverage_108,
  output        io_coverage_109,
  output        io_coverage_110,
  output        io_coverage_111,
  output        io_coverage_112,
  output        io_coverage_113,
  output        io_coverage_114,
  output        io_coverage_115,
  output        io_coverage_116,
  output        io_coverage_117,
  output        io_coverage_118,
  output        io_coverage_119,
  output        io_coverage_120,
  output        io_coverage_121,
  output        io_coverage_122,
  output        io_coverage_123,
  output        io_coverage_124,
  output        io_coverage_125,
  output        io_coverage_126,
  output        io_coverage_127,
  output        io_coverage_128,
  output        io_coverage_129,
  output        io_coverage_130,
  output        io_coverage_131,
  output        io_coverage_132,
  output        io_coverage_133,
  output        io_coverage_134,
  output        io_coverage_135,
  output        io_coverage_136,
  output        io_coverage_137,
  output        io_coverage_138,
  output        io_coverage_139,
  output        io_coverage_140,
  output        io_coverage_141,
  output        io_coverage_142,
  output        io_coverage_143,
  output        io_coverage_144,
  output        io_coverage_145,
  output        io_coverage_146,
  output        io_coverage_147,
  output        io_coverage_148,
  output        io_coverage_149,
  output        io_coverage_150,
  output        io_coverage_151,
  output        io_coverage_152,
  output        io_coverage_153,
  output        io_coverage_154,
  output        io_coverage_155,
  output        io_coverage_156,
  output        io_coverage_157,
  output        io_coverage_158,
  output        io_coverage_159,
  output        io_coverage_160,
  output        io_coverage_161,
  output        io_coverage_162,
  output        io_coverage_163,
  output        io_coverage_164,
  output        io_coverage_165,
  output        io_coverage_166,
  output        io_coverage_167,
  output        io_coverage_168,
  output        io_coverage_169,
  output        io_coverage_170,
  output        io_coverage_171,
  output        io_coverage_172,
  output        io_coverage_173,
  output        io_coverage_174,
  output        io_coverage_175,
  output        io_coverage_176,
  output        io_coverage_177,
  output        io_coverage_178,
  output        io_coverage_179,
  output        io_coverage_180,
  output        io_coverage_181,
  output        io_coverage_182,
  output        io_coverage_183,
  output        io_coverage_184,
  output        io_coverage_185,
  output        io_coverage_186
);
  wire [615:0] bb_auto_cover_out; // @[DUT.scala 29:24]
  wire  bb_assert_out; // @[DUT.scala 29:24]
  wire  bb_io_reset; // @[DUT.scala 29:24]
  wire  bb_io_imem_resp_valid; // @[DUT.scala 29:24]
  wire  bb_io_imem_req_ready; // @[DUT.scala 29:24]
  wire [31:0] bb_io_imem_resp_bits_data; // @[DUT.scala 29:24]
  wire  bb_metaReset; // @[DUT.scala 29:24]
  wire  bb_reset; // @[DUT.scala 29:24]
  wire  bb_clock; // @[DUT.scala 29:24]
  Sodor3Stage bb ( // @[DUT.scala 29:24]
    .auto_cover_out(bb_auto_cover_out),
    .assert_out(bb_assert_out),
    .io_reset(bb_io_reset),
    .io_imem_resp_valid(bb_io_imem_resp_valid),
    .io_imem_req_ready(bb_io_imem_req_ready),
    .io_imem_resp_bits_data(bb_io_imem_resp_bits_data),
    .metaReset(bb_metaReset),
    .reset(bb_reset),
    .clock(bb_clock)
  );
  assign io_coverage_0 = bb_assert_out; // @[DUT.scala 51:33]
  assign io_coverage_1 = bb_auto_cover_out[615]; // @[DUT.scala 51:33]
  assign io_coverage_2 = bb_auto_cover_out[614]; // @[DUT.scala 51:33]
  assign io_coverage_3 = bb_auto_cover_out[605]; // @[DUT.scala 51:33]
  assign io_coverage_4 = bb_auto_cover_out[604]; // @[DUT.scala 51:33]
  assign io_coverage_5 = bb_auto_cover_out[603]; // @[DUT.scala 51:33]
  assign io_coverage_6 = bb_auto_cover_out[602]; // @[DUT.scala 51:33]
  assign io_coverage_7 = bb_auto_cover_out[601]; // @[DUT.scala 51:33]
  assign io_coverage_8 = bb_auto_cover_out[600]; // @[DUT.scala 51:33]
  assign io_coverage_9 = bb_auto_cover_out[599]; // @[DUT.scala 51:33]
  assign io_coverage_10 = bb_auto_cover_out[598]; // @[DUT.scala 51:33]
  assign io_coverage_11 = bb_auto_cover_out[597]; // @[DUT.scala 51:33]
  assign io_coverage_12 = bb_auto_cover_out[596]; // @[DUT.scala 51:33]
  assign io_coverage_13 = bb_auto_cover_out[595]; // @[DUT.scala 51:33]
  assign io_coverage_14 = bb_auto_cover_out[594]; // @[DUT.scala 51:33]
  assign io_coverage_15 = bb_auto_cover_out[593]; // @[DUT.scala 51:33]
  assign io_coverage_16 = bb_auto_cover_out[592]; // @[DUT.scala 51:33]
  assign io_coverage_17 = bb_auto_cover_out[591]; // @[DUT.scala 51:33]
  assign io_coverage_18 = bb_auto_cover_out[590]; // @[DUT.scala 51:33]
  assign io_coverage_19 = bb_auto_cover_out[589]; // @[DUT.scala 51:33]
  assign io_coverage_20 = bb_auto_cover_out[588]; // @[DUT.scala 51:33]
  assign io_coverage_21 = bb_auto_cover_out[587]; // @[DUT.scala 51:33]
  assign io_coverage_22 = bb_auto_cover_out[586]; // @[DUT.scala 51:33]
  assign io_coverage_23 = bb_auto_cover_out[585]; // @[DUT.scala 51:33]
  assign io_coverage_24 = bb_auto_cover_out[584]; // @[DUT.scala 51:33]
  assign io_coverage_25 = bb_auto_cover_out[583]; // @[DUT.scala 51:33]
  assign io_coverage_26 = bb_auto_cover_out[582]; // @[DUT.scala 51:33]
  assign io_coverage_27 = bb_auto_cover_out[581]; // @[DUT.scala 51:33]
  assign io_coverage_28 = bb_auto_cover_out[580]; // @[DUT.scala 51:33]
  assign io_coverage_29 = bb_auto_cover_out[579]; // @[DUT.scala 51:33]
  assign io_coverage_30 = bb_auto_cover_out[578]; // @[DUT.scala 51:33]
  assign io_coverage_31 = bb_auto_cover_out[577]; // @[DUT.scala 51:33]
  assign io_coverage_32 = bb_auto_cover_out[576]; // @[DUT.scala 51:33]
  assign io_coverage_33 = bb_auto_cover_out[575]; // @[DUT.scala 51:33]
  assign io_coverage_34 = bb_auto_cover_out[574]; // @[DUT.scala 51:33]
  assign io_coverage_35 = bb_auto_cover_out[573]; // @[DUT.scala 51:33]
  assign io_coverage_36 = bb_auto_cover_out[572]; // @[DUT.scala 51:33]
  assign io_coverage_37 = bb_auto_cover_out[571]; // @[DUT.scala 51:33]
  assign io_coverage_38 = bb_auto_cover_out[570]; // @[DUT.scala 51:33]
  assign io_coverage_39 = bb_auto_cover_out[569]; // @[DUT.scala 51:33]
  assign io_coverage_40 = bb_auto_cover_out[540]; // @[DUT.scala 51:33]
  assign io_coverage_41 = bb_auto_cover_out[539]; // @[DUT.scala 51:33]
  assign io_coverage_42 = bb_auto_cover_out[538]; // @[DUT.scala 51:33]
  assign io_coverage_43 = bb_auto_cover_out[537]; // @[DUT.scala 51:33]
  assign io_coverage_44 = bb_auto_cover_out[536]; // @[DUT.scala 51:33]
  assign io_coverage_45 = bb_auto_cover_out[535]; // @[DUT.scala 51:33]
  assign io_coverage_46 = bb_auto_cover_out[357]; // @[DUT.scala 51:33]
  assign io_coverage_47 = bb_auto_cover_out[356]; // @[DUT.scala 51:33]
  assign io_coverage_48 = bb_auto_cover_out[355]; // @[DUT.scala 51:33]
  assign io_coverage_49 = bb_auto_cover_out[354]; // @[DUT.scala 51:33]
  assign io_coverage_50 = bb_auto_cover_out[353]; // @[DUT.scala 51:33]
  assign io_coverage_51 = bb_auto_cover_out[309]; // @[DUT.scala 51:33]
  assign io_coverage_52 = bb_auto_cover_out[308]; // @[DUT.scala 51:33]
  assign io_coverage_53 = bb_auto_cover_out[307]; // @[DUT.scala 51:33]
  assign io_coverage_54 = bb_auto_cover_out[306]; // @[DUT.scala 51:33]
  assign io_coverage_55 = bb_auto_cover_out[305]; // @[DUT.scala 51:33]
  assign io_coverage_56 = bb_auto_cover_out[304]; // @[DUT.scala 51:33]
  assign io_coverage_57 = bb_auto_cover_out[303]; // @[DUT.scala 51:33]
  assign io_coverage_58 = bb_auto_cover_out[302]; // @[DUT.scala 51:33]
  assign io_coverage_59 = bb_auto_cover_out[301]; // @[DUT.scala 51:33]
  assign io_coverage_60 = bb_auto_cover_out[300]; // @[DUT.scala 51:33]
  assign io_coverage_61 = bb_auto_cover_out[299]; // @[DUT.scala 51:33]
  assign io_coverage_62 = bb_auto_cover_out[298]; // @[DUT.scala 51:33]
  assign io_coverage_63 = bb_auto_cover_out[297]; // @[DUT.scala 51:33]
  assign io_coverage_64 = bb_auto_cover_out[296]; // @[DUT.scala 51:33]
  assign io_coverage_65 = bb_auto_cover_out[295]; // @[DUT.scala 51:33]
  assign io_coverage_66 = bb_auto_cover_out[294]; // @[DUT.scala 51:33]
  assign io_coverage_67 = bb_auto_cover_out[293]; // @[DUT.scala 51:33]
  assign io_coverage_68 = bb_auto_cover_out[286]; // @[DUT.scala 51:33]
  assign io_coverage_69 = bb_auto_cover_out[281]; // @[DUT.scala 51:33]
  assign io_coverage_70 = bb_auto_cover_out[280]; // @[DUT.scala 51:33]
  assign io_coverage_71 = bb_auto_cover_out[279]; // @[DUT.scala 51:33]
  assign io_coverage_72 = bb_auto_cover_out[278]; // @[DUT.scala 51:33]
  assign io_coverage_73 = bb_auto_cover_out[277]; // @[DUT.scala 51:33]
  assign io_coverage_74 = bb_auto_cover_out[276]; // @[DUT.scala 51:33]
  assign io_coverage_75 = bb_auto_cover_out[275]; // @[DUT.scala 51:33]
  assign io_coverage_76 = bb_auto_cover_out[274]; // @[DUT.scala 51:33]
  assign io_coverage_77 = bb_auto_cover_out[272]; // @[DUT.scala 51:33]
  assign io_coverage_78 = bb_auto_cover_out[271]; // @[DUT.scala 51:33]
  assign io_coverage_79 = bb_auto_cover_out[268]; // @[DUT.scala 51:33]
  assign io_coverage_80 = bb_auto_cover_out[267]; // @[DUT.scala 51:33]
  assign io_coverage_81 = bb_auto_cover_out[266]; // @[DUT.scala 51:33]
  assign io_coverage_82 = bb_auto_cover_out[263]; // @[DUT.scala 51:33]
  assign io_coverage_83 = bb_auto_cover_out[261]; // @[DUT.scala 51:33]
  assign io_coverage_84 = bb_auto_cover_out[259]; // @[DUT.scala 51:33]
  assign io_coverage_85 = bb_auto_cover_out[258]; // @[DUT.scala 51:33]
  assign io_coverage_86 = bb_auto_cover_out[257]; // @[DUT.scala 51:33]
  assign io_coverage_87 = bb_auto_cover_out[256]; // @[DUT.scala 51:33]
  assign io_coverage_88 = bb_auto_cover_out[255]; // @[DUT.scala 51:33]
  assign io_coverage_89 = bb_auto_cover_out[254]; // @[DUT.scala 51:33]
  assign io_coverage_90 = bb_auto_cover_out[253]; // @[DUT.scala 51:33]
  assign io_coverage_91 = bb_auto_cover_out[252]; // @[DUT.scala 51:33]
  assign io_coverage_92 = bb_auto_cover_out[251]; // @[DUT.scala 51:33]
  assign io_coverage_93 = bb_auto_cover_out[250]; // @[DUT.scala 51:33]
  assign io_coverage_94 = bb_auto_cover_out[249]; // @[DUT.scala 51:33]
  assign io_coverage_95 = bb_auto_cover_out[248]; // @[DUT.scala 51:33]
  assign io_coverage_96 = bb_auto_cover_out[247]; // @[DUT.scala 51:33]
  assign io_coverage_97 = bb_auto_cover_out[246]; // @[DUT.scala 51:33]
  assign io_coverage_98 = bb_auto_cover_out[245]; // @[DUT.scala 51:33]
  assign io_coverage_99 = bb_auto_cover_out[244]; // @[DUT.scala 51:33]
  assign io_coverage_100 = bb_auto_cover_out[243]; // @[DUT.scala 51:33]
  assign io_coverage_101 = bb_auto_cover_out[242]; // @[DUT.scala 51:33]
  assign io_coverage_102 = bb_auto_cover_out[241]; // @[DUT.scala 51:33]
  assign io_coverage_103 = bb_auto_cover_out[240]; // @[DUT.scala 51:33]
  assign io_coverage_104 = bb_auto_cover_out[239]; // @[DUT.scala 51:33]
  assign io_coverage_105 = bb_auto_cover_out[238]; // @[DUT.scala 51:33]
  assign io_coverage_106 = bb_auto_cover_out[237]; // @[DUT.scala 51:33]
  assign io_coverage_107 = bb_auto_cover_out[236]; // @[DUT.scala 51:33]
  assign io_coverage_108 = bb_auto_cover_out[235]; // @[DUT.scala 51:33]
  assign io_coverage_109 = bb_auto_cover_out[234]; // @[DUT.scala 51:33]
  assign io_coverage_110 = bb_auto_cover_out[233]; // @[DUT.scala 51:33]
  assign io_coverage_111 = bb_auto_cover_out[232]; // @[DUT.scala 51:33]
  assign io_coverage_112 = bb_auto_cover_out[231]; // @[DUT.scala 51:33]
  assign io_coverage_113 = bb_auto_cover_out[230]; // @[DUT.scala 51:33]
  assign io_coverage_114 = bb_auto_cover_out[229]; // @[DUT.scala 51:33]
  assign io_coverage_115 = bb_auto_cover_out[228]; // @[DUT.scala 51:33]
  assign io_coverage_116 = bb_auto_cover_out[227]; // @[DUT.scala 51:33]
  assign io_coverage_117 = bb_auto_cover_out[226]; // @[DUT.scala 51:33]
  assign io_coverage_118 = bb_auto_cover_out[225]; // @[DUT.scala 51:33]
  assign io_coverage_119 = bb_auto_cover_out[224]; // @[DUT.scala 51:33]
  assign io_coverage_120 = bb_auto_cover_out[223]; // @[DUT.scala 51:33]
  assign io_coverage_121 = bb_auto_cover_out[222]; // @[DUT.scala 51:33]
  assign io_coverage_122 = bb_auto_cover_out[221]; // @[DUT.scala 51:33]
  assign io_coverage_123 = bb_auto_cover_out[220]; // @[DUT.scala 51:33]
  assign io_coverage_124 = bb_auto_cover_out[219]; // @[DUT.scala 51:33]
  assign io_coverage_125 = bb_auto_cover_out[218]; // @[DUT.scala 51:33]
  assign io_coverage_126 = bb_auto_cover_out[217]; // @[DUT.scala 51:33]
  assign io_coverage_127 = bb_auto_cover_out[216]; // @[DUT.scala 51:33]
  assign io_coverage_128 = bb_auto_cover_out[215]; // @[DUT.scala 51:33]
  assign io_coverage_129 = bb_auto_cover_out[214]; // @[DUT.scala 51:33]
  assign io_coverage_130 = bb_auto_cover_out[213]; // @[DUT.scala 51:33]
  assign io_coverage_131 = bb_auto_cover_out[212]; // @[DUT.scala 51:33]
  assign io_coverage_132 = bb_auto_cover_out[211]; // @[DUT.scala 51:33]
  assign io_coverage_133 = bb_auto_cover_out[210]; // @[DUT.scala 51:33]
  assign io_coverage_134 = bb_auto_cover_out[209]; // @[DUT.scala 51:33]
  assign io_coverage_135 = bb_auto_cover_out[208]; // @[DUT.scala 51:33]
  assign io_coverage_136 = bb_auto_cover_out[207]; // @[DUT.scala 51:33]
  assign io_coverage_137 = bb_auto_cover_out[206]; // @[DUT.scala 51:33]
  assign io_coverage_138 = bb_auto_cover_out[205]; // @[DUT.scala 51:33]
  assign io_coverage_139 = bb_auto_cover_out[204]; // @[DUT.scala 51:33]
  assign io_coverage_140 = bb_auto_cover_out[203]; // @[DUT.scala 51:33]
  assign io_coverage_141 = bb_auto_cover_out[202]; // @[DUT.scala 51:33]
  assign io_coverage_142 = bb_auto_cover_out[201]; // @[DUT.scala 51:33]
  assign io_coverage_143 = bb_auto_cover_out[200]; // @[DUT.scala 51:33]
  assign io_coverage_144 = bb_auto_cover_out[199]; // @[DUT.scala 51:33]
  assign io_coverage_145 = bb_auto_cover_out[198]; // @[DUT.scala 51:33]
  assign io_coverage_146 = bb_auto_cover_out[197]; // @[DUT.scala 51:33]
  assign io_coverage_147 = bb_auto_cover_out[196]; // @[DUT.scala 51:33]
  assign io_coverage_148 = bb_auto_cover_out[195]; // @[DUT.scala 51:33]
  assign io_coverage_149 = bb_auto_cover_out[194]; // @[DUT.scala 51:33]
  assign io_coverage_150 = bb_auto_cover_out[193]; // @[DUT.scala 51:33]
  assign io_coverage_151 = bb_auto_cover_out[192]; // @[DUT.scala 51:33]
  assign io_coverage_152 = bb_auto_cover_out[191]; // @[DUT.scala 51:33]
  assign io_coverage_153 = bb_auto_cover_out[190]; // @[DUT.scala 51:33]
  assign io_coverage_154 = bb_auto_cover_out[189]; // @[DUT.scala 51:33]
  assign io_coverage_155 = bb_auto_cover_out[188]; // @[DUT.scala 51:33]
  assign io_coverage_156 = bb_auto_cover_out[187]; // @[DUT.scala 51:33]
  assign io_coverage_157 = bb_auto_cover_out[186]; // @[DUT.scala 51:33]
  assign io_coverage_158 = bb_auto_cover_out[185]; // @[DUT.scala 51:33]
  assign io_coverage_159 = bb_auto_cover_out[184]; // @[DUT.scala 51:33]
  assign io_coverage_160 = bb_auto_cover_out[183]; // @[DUT.scala 51:33]
  assign io_coverage_161 = bb_auto_cover_out[182]; // @[DUT.scala 51:33]
  assign io_coverage_162 = bb_auto_cover_out[181]; // @[DUT.scala 51:33]
  assign io_coverage_163 = bb_auto_cover_out[180]; // @[DUT.scala 51:33]
  assign io_coverage_164 = bb_auto_cover_out[179]; // @[DUT.scala 51:33]
  assign io_coverage_165 = bb_auto_cover_out[107]; // @[DUT.scala 51:33]
  assign io_coverage_166 = bb_auto_cover_out[103]; // @[DUT.scala 51:33]
  assign io_coverage_167 = bb_auto_cover_out[92]; // @[DUT.scala 51:33]
  assign io_coverage_168 = bb_auto_cover_out[29]; // @[DUT.scala 51:33]
  assign io_coverage_169 = bb_auto_cover_out[28]; // @[DUT.scala 51:33]
  assign io_coverage_170 = bb_auto_cover_out[27]; // @[DUT.scala 51:33]
  assign io_coverage_171 = bb_auto_cover_out[26]; // @[DUT.scala 51:33]
  assign io_coverage_172 = bb_auto_cover_out[25]; // @[DUT.scala 51:33]
  assign io_coverage_173 = bb_auto_cover_out[24]; // @[DUT.scala 51:33]
  assign io_coverage_174 = bb_auto_cover_out[23]; // @[DUT.scala 51:33]
  assign io_coverage_175 = bb_auto_cover_out[22]; // @[DUT.scala 51:33]
  assign io_coverage_176 = bb_auto_cover_out[21]; // @[DUT.scala 51:33]
  assign io_coverage_177 = bb_auto_cover_out[20]; // @[DUT.scala 51:33]
  assign io_coverage_178 = bb_auto_cover_out[19]; // @[DUT.scala 51:33]
  assign io_coverage_179 = bb_auto_cover_out[18]; // @[DUT.scala 51:33]
  assign io_coverage_180 = bb_auto_cover_out[16]; // @[DUT.scala 51:33]
  assign io_coverage_181 = bb_auto_cover_out[15]; // @[DUT.scala 51:33]
  assign io_coverage_182 = bb_auto_cover_out[14]; // @[DUT.scala 51:33]
  assign io_coverage_183 = bb_auto_cover_out[11]; // @[DUT.scala 51:33]
  assign io_coverage_184 = bb_auto_cover_out[9]; // @[DUT.scala 51:33]
  assign io_coverage_185 = bb_auto_cover_out[5]; // @[DUT.scala 51:33]
  assign io_coverage_186 = bb_auto_cover_out[4]; // @[DUT.scala 51:33]
  assign bb_io_reset = io_inputs[0]; // @[DUT.scala 40:25]
  assign bb_io_imem_resp_valid = io_inputs[1]; // @[DUT.scala 40:25]
  assign bb_io_imem_req_ready = io_inputs[2]; // @[DUT.scala 40:25]
  assign bb_io_imem_resp_bits_data = io_inputs[34:3]; // @[DUT.scala 40:25]
  assign bb_metaReset = io_meta_reset; // @[DUT.scala 35:27]
  assign bb_reset = reset; // @[DUT.scala 34:23]
  assign bb_clock = clock; // @[DUT.scala 33:23]
endmodule
module SaturatingCounter(
  input   clock,
  input   reset,
  input   io_enable,
  output  io_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  count; // @[coverage.scala 11:28]
  wire  _T = ~io_enable; // @[coverage.scala 14:22]
  wire  _T_2 = _T | count; // @[coverage.scala 14:33]
  wire  _T_4 = count + 1'h1; // @[coverage.scala 14:64]
  assign io_value = count; // @[coverage.scala 12:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      count <= 1'h0;
    end else if (!(_T_2)) begin
      count <= _T_4;
    end
  end
endmodule
module VerilatorHarness(
  input        clock,
  input        reset,
  input  [7:0] io_input_bytes_0,
  input  [7:0] io_input_bytes_1,
  input  [7:0] io_input_bytes_2,
  input  [7:0] io_input_bytes_3,
  input  [7:0] io_input_bytes_4,
  input  [7:0] io_input_bytes_5,
  input  [7:0] io_input_bytes_6,
  input  [7:0] io_input_bytes_7,
  output [7:0] io_coverage_bytes_0,
  output [7:0] io_coverage_bytes_1,
  output [7:0] io_coverage_bytes_2,
  output [7:0] io_coverage_bytes_3,
  output [7:0] io_coverage_bytes_4,
  output [7:0] io_coverage_bytes_5,
  output [7:0] io_coverage_bytes_6,
  output [7:0] io_coverage_bytes_7,
  output [7:0] io_coverage_bytes_8,
  output [7:0] io_coverage_bytes_9,
  output [7:0] io_coverage_bytes_10,
  output [7:0] io_coverage_bytes_11,
  output [7:0] io_coverage_bytes_12,
  output [7:0] io_coverage_bytes_13,
  output [7:0] io_coverage_bytes_14,
  output [7:0] io_coverage_bytes_15,
  output [7:0] io_coverage_bytes_16,
  output [7:0] io_coverage_bytes_17,
  output [7:0] io_coverage_bytes_18,
  output [7:0] io_coverage_bytes_19,
  output [7:0] io_coverage_bytes_20,
  output [7:0] io_coverage_bytes_21,
  output [7:0] io_coverage_bytes_22,
  output [7:0] io_coverage_bytes_23,
  output [7:0] io_coverage_bytes_24,
  output [7:0] io_coverage_bytes_25,
  output [7:0] io_coverage_bytes_26,
  output [7:0] io_coverage_bytes_27,
  output [7:0] io_coverage_bytes_28,
  output [7:0] io_coverage_bytes_29,
  output [7:0] io_coverage_bytes_30,
  output [7:0] io_coverage_bytes_31,
  output [7:0] io_coverage_bytes_32,
  output [7:0] io_coverage_bytes_33,
  output [7:0] io_coverage_bytes_34,
  output [7:0] io_coverage_bytes_35,
  output [7:0] io_coverage_bytes_36,
  output [7:0] io_coverage_bytes_37,
  output [7:0] io_coverage_bytes_38,
  output [7:0] io_coverage_bytes_39,
  output [7:0] io_coverage_bytes_40,
  output [7:0] io_coverage_bytes_41,
  output [7:0] io_coverage_bytes_42,
  output [7:0] io_coverage_bytes_43,
  output [7:0] io_coverage_bytes_44,
  output [7:0] io_coverage_bytes_45,
  output [7:0] io_coverage_bytes_46,
  output [7:0] io_coverage_bytes_47,
  output [7:0] io_coverage_bytes_48,
  output [7:0] io_coverage_bytes_49,
  output [7:0] io_coverage_bytes_50,
  output [7:0] io_coverage_bytes_51,
  output [7:0] io_coverage_bytes_52,
  output [7:0] io_coverage_bytes_53,
  output [7:0] io_coverage_bytes_54,
  output [7:0] io_coverage_bytes_55,
  output [7:0] io_coverage_bytes_56,
  output [7:0] io_coverage_bytes_57,
  output [7:0] io_coverage_bytes_58,
  output [7:0] io_coverage_bytes_59,
  output [7:0] io_coverage_bytes_60,
  output [7:0] io_coverage_bytes_61,
  output [7:0] io_coverage_bytes_62,
  output [7:0] io_coverage_bytes_63,
  output [7:0] io_coverage_bytes_64,
  output [7:0] io_coverage_bytes_65,
  output [7:0] io_coverage_bytes_66,
  output [7:0] io_coverage_bytes_67,
  output [7:0] io_coverage_bytes_68,
  output [7:0] io_coverage_bytes_69,
  output [7:0] io_coverage_bytes_70,
  output [7:0] io_coverage_bytes_71,
  output [7:0] io_coverage_bytes_72,
  output [7:0] io_coverage_bytes_73,
  output [7:0] io_coverage_bytes_74,
  output [7:0] io_coverage_bytes_75,
  output [7:0] io_coverage_bytes_76,
  output [7:0] io_coverage_bytes_77,
  output [7:0] io_coverage_bytes_78,
  output [7:0] io_coverage_bytes_79,
  output [7:0] io_coverage_bytes_80,
  output [7:0] io_coverage_bytes_81,
  output [7:0] io_coverage_bytes_82,
  output [7:0] io_coverage_bytes_83,
  output [7:0] io_coverage_bytes_84,
  output [7:0] io_coverage_bytes_85,
  output [7:0] io_coverage_bytes_86,
  output [7:0] io_coverage_bytes_87,
  output [7:0] io_coverage_bytes_88,
  output [7:0] io_coverage_bytes_89,
  output [7:0] io_coverage_bytes_90,
  output [7:0] io_coverage_bytes_91,
  output [7:0] io_coverage_bytes_92,
  output [7:0] io_coverage_bytes_93,
  output [7:0] io_coverage_bytes_94,
  output [7:0] io_coverage_bytes_95,
  output [7:0] io_coverage_bytes_96,
  output [7:0] io_coverage_bytes_97,
  output [7:0] io_coverage_bytes_98,
  output [7:0] io_coverage_bytes_99,
  output [7:0] io_coverage_bytes_100,
  output [7:0] io_coverage_bytes_101,
  output [7:0] io_coverage_bytes_102,
  output [7:0] io_coverage_bytes_103,
  output [7:0] io_coverage_bytes_104,
  output [7:0] io_coverage_bytes_105,
  output [7:0] io_coverage_bytes_106,
  output [7:0] io_coverage_bytes_107,
  output [7:0] io_coverage_bytes_108,
  output [7:0] io_coverage_bytes_109,
  output [7:0] io_coverage_bytes_110,
  output [7:0] io_coverage_bytes_111,
  output [7:0] io_coverage_bytes_112,
  output [7:0] io_coverage_bytes_113,
  output [7:0] io_coverage_bytes_114,
  output [7:0] io_coverage_bytes_115,
  output [7:0] io_coverage_bytes_116,
  output [7:0] io_coverage_bytes_117,
  output [7:0] io_coverage_bytes_118,
  output [7:0] io_coverage_bytes_119,
  output [7:0] io_coverage_bytes_120,
  output [7:0] io_coverage_bytes_121,
  output [7:0] io_coverage_bytes_122,
  output [7:0] io_coverage_bytes_123,
  output [7:0] io_coverage_bytes_124,
  output [7:0] io_coverage_bytes_125,
  output [7:0] io_coverage_bytes_126,
  output [7:0] io_coverage_bytes_127,
  output [7:0] io_coverage_bytes_128,
  output [7:0] io_coverage_bytes_129,
  output [7:0] io_coverage_bytes_130,
  output [7:0] io_coverage_bytes_131,
  output [7:0] io_coverage_bytes_132,
  output [7:0] io_coverage_bytes_133,
  output [7:0] io_coverage_bytes_134,
  output [7:0] io_coverage_bytes_135,
  output [7:0] io_coverage_bytes_136,
  output [7:0] io_coverage_bytes_137,
  output [7:0] io_coverage_bytes_138,
  output [7:0] io_coverage_bytes_139,
  output [7:0] io_coverage_bytes_140,
  output [7:0] io_coverage_bytes_141,
  output [7:0] io_coverage_bytes_142,
  output [7:0] io_coverage_bytes_143,
  output [7:0] io_coverage_bytes_144,
  output [7:0] io_coverage_bytes_145,
  output [7:0] io_coverage_bytes_146,
  output [7:0] io_coverage_bytes_147,
  output [7:0] io_coverage_bytes_148,
  output [7:0] io_coverage_bytes_149,
  output [7:0] io_coverage_bytes_150,
  output [7:0] io_coverage_bytes_151,
  output [7:0] io_coverage_bytes_152,
  output [7:0] io_coverage_bytes_153,
  output [7:0] io_coverage_bytes_154,
  output [7:0] io_coverage_bytes_155,
  output [7:0] io_coverage_bytes_156,
  output [7:0] io_coverage_bytes_157,
  output [7:0] io_coverage_bytes_158,
  output [7:0] io_coverage_bytes_159,
  output [7:0] io_coverage_bytes_160,
  output [7:0] io_coverage_bytes_161,
  output [7:0] io_coverage_bytes_162,
  output [7:0] io_coverage_bytes_163,
  output [7:0] io_coverage_bytes_164,
  output [7:0] io_coverage_bytes_165,
  output [7:0] io_coverage_bytes_166,
  output [7:0] io_coverage_bytes_167,
  output [7:0] io_coverage_bytes_168,
  output [7:0] io_coverage_bytes_169,
  output [7:0] io_coverage_bytes_170,
  output [7:0] io_coverage_bytes_171,
  output [7:0] io_coverage_bytes_172,
  output [7:0] io_coverage_bytes_173,
  output [7:0] io_coverage_bytes_174,
  output [7:0] io_coverage_bytes_175,
  output [7:0] io_coverage_bytes_176,
  output [7:0] io_coverage_bytes_177,
  output [7:0] io_coverage_bytes_178,
  output [7:0] io_coverage_bytes_179,
  output [7:0] io_coverage_bytes_180,
  output [7:0] io_coverage_bytes_181,
  output [7:0] io_coverage_bytes_182,
  output [7:0] io_coverage_bytes_183,
  output [7:0] io_coverage_bytes_184,
  output [7:0] io_coverage_bytes_185,
  output [7:0] io_coverage_bytes_186,
  output [7:0] io_coverage_bytes_187,
  output [7:0] io_coverage_bytes_188,
  output [7:0] io_coverage_bytes_189,
  input        io_meta_reset
);
  wire  dut_clock; // @[VerilatorHarness.scala 42:25]
  wire  dut_reset; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_meta_reset; // @[VerilatorHarness.scala 42:25]
  wire [34:0] dut_io_inputs; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_0; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_1; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_2; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_3; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_4; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_5; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_6; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_7; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_8; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_9; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_10; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_11; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_12; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_13; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_14; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_15; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_16; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_17; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_18; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_19; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_20; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_21; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_22; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_23; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_24; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_25; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_26; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_27; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_28; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_29; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_30; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_31; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_32; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_33; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_34; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_35; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_36; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_37; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_38; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_39; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_40; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_41; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_42; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_43; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_44; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_45; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_46; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_47; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_48; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_49; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_50; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_51; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_52; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_53; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_54; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_55; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_56; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_57; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_58; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_59; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_60; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_61; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_62; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_63; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_64; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_65; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_66; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_67; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_68; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_69; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_70; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_71; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_72; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_73; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_74; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_75; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_76; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_77; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_78; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_79; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_80; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_81; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_82; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_83; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_84; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_85; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_86; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_87; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_88; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_89; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_90; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_91; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_92; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_93; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_94; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_95; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_96; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_97; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_98; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_99; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_100; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_101; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_102; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_103; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_104; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_105; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_106; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_107; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_108; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_109; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_110; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_111; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_112; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_113; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_114; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_115; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_116; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_117; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_118; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_119; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_120; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_121; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_122; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_123; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_124; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_125; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_126; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_127; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_128; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_129; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_130; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_131; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_132; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_133; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_134; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_135; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_136; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_137; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_138; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_139; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_140; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_141; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_142; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_143; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_144; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_145; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_146; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_147; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_148; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_149; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_150; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_151; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_152; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_153; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_154; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_155; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_156; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_157; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_158; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_159; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_160; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_161; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_162; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_163; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_164; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_165; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_166; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_167; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_168; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_169; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_170; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_171; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_172; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_173; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_174; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_175; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_176; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_177; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_178; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_179; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_180; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_181; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_182; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_183; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_184; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_185; // @[VerilatorHarness.scala 42:25]
  wire  dut_io_coverage_186; // @[VerilatorHarness.scala 42:25]
  wire  SaturatingCounter_clock; // @[coverage.scala 121:35]
  wire  SaturatingCounter_reset; // @[coverage.scala 121:35]
  wire  SaturatingCounter_io_enable; // @[coverage.scala 121:35]
  wire  SaturatingCounter_io_value; // @[coverage.scala 121:35]
  wire  SaturatingCounter_1_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_1_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_1_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_1_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_2_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_2_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_2_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_2_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_3_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_3_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_3_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_3_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_4_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_4_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_4_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_4_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_5_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_5_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_5_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_5_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_6_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_6_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_6_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_6_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_7_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_7_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_7_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_7_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_8_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_8_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_8_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_8_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_9_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_9_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_9_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_9_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_10_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_10_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_10_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_10_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_11_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_11_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_11_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_11_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_12_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_12_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_12_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_12_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_13_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_13_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_13_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_13_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_14_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_14_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_14_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_14_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_15_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_15_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_15_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_15_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_16_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_16_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_16_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_16_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_17_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_17_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_17_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_17_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_18_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_18_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_18_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_18_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_19_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_19_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_19_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_19_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_20_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_20_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_20_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_20_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_21_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_21_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_21_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_21_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_22_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_22_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_22_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_22_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_23_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_23_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_23_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_23_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_24_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_24_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_24_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_24_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_25_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_25_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_25_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_25_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_26_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_26_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_26_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_26_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_27_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_27_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_27_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_27_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_28_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_28_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_28_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_28_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_29_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_29_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_29_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_29_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_30_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_30_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_30_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_30_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_31_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_31_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_31_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_31_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_32_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_32_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_32_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_32_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_33_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_33_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_33_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_33_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_34_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_34_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_34_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_34_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_35_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_35_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_35_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_35_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_36_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_36_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_36_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_36_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_37_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_37_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_37_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_37_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_38_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_38_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_38_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_38_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_39_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_39_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_39_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_39_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_40_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_40_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_40_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_40_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_41_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_41_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_41_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_41_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_42_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_42_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_42_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_42_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_43_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_43_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_43_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_43_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_44_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_44_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_44_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_44_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_45_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_45_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_45_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_45_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_46_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_46_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_46_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_46_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_47_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_47_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_47_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_47_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_48_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_48_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_48_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_48_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_49_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_49_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_49_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_49_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_50_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_50_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_50_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_50_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_51_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_51_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_51_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_51_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_52_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_52_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_52_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_52_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_53_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_53_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_53_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_53_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_54_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_54_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_54_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_54_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_55_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_55_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_55_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_55_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_56_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_56_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_56_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_56_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_57_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_57_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_57_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_57_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_58_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_58_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_58_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_58_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_59_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_59_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_59_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_59_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_60_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_60_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_60_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_60_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_61_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_61_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_61_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_61_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_62_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_62_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_62_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_62_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_63_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_63_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_63_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_63_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_64_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_64_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_64_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_64_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_65_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_65_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_65_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_65_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_66_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_66_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_66_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_66_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_67_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_67_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_67_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_67_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_68_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_68_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_68_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_68_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_69_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_69_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_69_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_69_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_70_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_70_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_70_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_70_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_71_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_71_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_71_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_71_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_72_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_72_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_72_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_72_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_73_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_73_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_73_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_73_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_74_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_74_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_74_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_74_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_75_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_75_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_75_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_75_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_76_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_76_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_76_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_76_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_77_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_77_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_77_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_77_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_78_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_78_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_78_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_78_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_79_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_79_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_79_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_79_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_80_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_80_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_80_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_80_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_81_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_81_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_81_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_81_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_82_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_82_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_82_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_82_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_83_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_83_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_83_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_83_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_84_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_84_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_84_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_84_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_85_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_85_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_85_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_85_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_86_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_86_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_86_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_86_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_87_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_87_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_87_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_87_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_88_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_88_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_88_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_88_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_89_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_89_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_89_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_89_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_90_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_90_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_90_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_90_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_91_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_91_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_91_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_91_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_92_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_92_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_92_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_92_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_93_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_93_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_93_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_93_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_94_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_94_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_94_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_94_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_95_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_95_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_95_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_95_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_96_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_96_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_96_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_96_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_97_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_97_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_97_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_97_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_98_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_98_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_98_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_98_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_99_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_99_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_99_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_99_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_100_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_100_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_100_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_100_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_101_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_101_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_101_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_101_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_102_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_102_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_102_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_102_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_103_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_103_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_103_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_103_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_104_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_104_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_104_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_104_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_105_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_105_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_105_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_105_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_106_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_106_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_106_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_106_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_107_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_107_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_107_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_107_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_108_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_108_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_108_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_108_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_109_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_109_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_109_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_109_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_110_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_110_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_110_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_110_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_111_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_111_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_111_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_111_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_112_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_112_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_112_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_112_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_113_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_113_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_113_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_113_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_114_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_114_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_114_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_114_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_115_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_115_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_115_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_115_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_116_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_116_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_116_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_116_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_117_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_117_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_117_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_117_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_118_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_118_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_118_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_118_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_119_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_119_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_119_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_119_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_120_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_120_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_120_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_120_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_121_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_121_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_121_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_121_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_122_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_122_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_122_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_122_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_123_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_123_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_123_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_123_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_124_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_124_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_124_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_124_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_125_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_125_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_125_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_125_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_126_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_126_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_126_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_126_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_127_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_127_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_127_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_127_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_128_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_128_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_128_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_128_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_129_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_129_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_129_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_129_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_130_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_130_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_130_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_130_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_131_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_131_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_131_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_131_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_132_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_132_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_132_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_132_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_133_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_133_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_133_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_133_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_134_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_134_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_134_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_134_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_135_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_135_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_135_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_135_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_136_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_136_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_136_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_136_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_137_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_137_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_137_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_137_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_138_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_138_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_138_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_138_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_139_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_139_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_139_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_139_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_140_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_140_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_140_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_140_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_141_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_141_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_141_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_141_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_142_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_142_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_142_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_142_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_143_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_143_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_143_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_143_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_144_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_144_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_144_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_144_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_145_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_145_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_145_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_145_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_146_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_146_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_146_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_146_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_147_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_147_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_147_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_147_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_148_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_148_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_148_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_148_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_149_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_149_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_149_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_149_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_150_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_150_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_150_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_150_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_151_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_151_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_151_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_151_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_152_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_152_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_152_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_152_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_153_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_153_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_153_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_153_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_154_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_154_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_154_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_154_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_155_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_155_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_155_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_155_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_156_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_156_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_156_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_156_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_157_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_157_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_157_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_157_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_158_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_158_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_158_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_158_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_159_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_159_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_159_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_159_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_160_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_160_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_160_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_160_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_161_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_161_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_161_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_161_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_162_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_162_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_162_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_162_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_163_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_163_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_163_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_163_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_164_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_164_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_164_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_164_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_165_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_165_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_165_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_165_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_166_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_166_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_166_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_166_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_167_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_167_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_167_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_167_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_168_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_168_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_168_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_168_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_169_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_169_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_169_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_169_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_170_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_170_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_170_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_170_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_171_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_171_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_171_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_171_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_172_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_172_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_172_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_172_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_173_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_173_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_173_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_173_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_174_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_174_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_174_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_174_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_175_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_175_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_175_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_175_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_176_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_176_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_176_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_176_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_177_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_177_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_177_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_177_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_178_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_178_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_178_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_178_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_179_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_179_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_179_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_179_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_180_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_180_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_180_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_180_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_181_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_181_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_181_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_181_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_182_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_182_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_182_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_182_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_183_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_183_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_183_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_183_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_184_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_184_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_184_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_184_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_185_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_185_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_185_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_185_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_186_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_186_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_186_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_186_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_187_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_187_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_187_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_187_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_188_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_188_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_188_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_188_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_189_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_189_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_189_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_189_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_190_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_190_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_190_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_190_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_191_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_191_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_191_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_191_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_192_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_192_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_192_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_192_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_193_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_193_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_193_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_193_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_194_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_194_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_194_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_194_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_195_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_195_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_195_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_195_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_196_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_196_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_196_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_196_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_197_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_197_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_197_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_197_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_198_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_198_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_198_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_198_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_199_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_199_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_199_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_199_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_200_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_200_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_200_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_200_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_201_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_201_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_201_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_201_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_202_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_202_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_202_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_202_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_203_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_203_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_203_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_203_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_204_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_204_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_204_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_204_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_205_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_205_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_205_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_205_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_206_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_206_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_206_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_206_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_207_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_207_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_207_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_207_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_208_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_208_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_208_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_208_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_209_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_209_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_209_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_209_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_210_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_210_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_210_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_210_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_211_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_211_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_211_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_211_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_212_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_212_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_212_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_212_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_213_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_213_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_213_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_213_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_214_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_214_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_214_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_214_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_215_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_215_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_215_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_215_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_216_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_216_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_216_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_216_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_217_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_217_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_217_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_217_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_218_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_218_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_218_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_218_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_219_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_219_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_219_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_219_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_220_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_220_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_220_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_220_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_221_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_221_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_221_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_221_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_222_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_222_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_222_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_222_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_223_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_223_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_223_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_223_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_224_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_224_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_224_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_224_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_225_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_225_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_225_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_225_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_226_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_226_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_226_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_226_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_227_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_227_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_227_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_227_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_228_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_228_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_228_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_228_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_229_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_229_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_229_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_229_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_230_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_230_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_230_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_230_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_231_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_231_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_231_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_231_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_232_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_232_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_232_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_232_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_233_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_233_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_233_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_233_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_234_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_234_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_234_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_234_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_235_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_235_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_235_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_235_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_236_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_236_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_236_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_236_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_237_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_237_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_237_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_237_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_238_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_238_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_238_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_238_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_239_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_239_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_239_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_239_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_240_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_240_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_240_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_240_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_241_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_241_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_241_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_241_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_242_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_242_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_242_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_242_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_243_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_243_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_243_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_243_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_244_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_244_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_244_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_244_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_245_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_245_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_245_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_245_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_246_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_246_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_246_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_246_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_247_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_247_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_247_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_247_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_248_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_248_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_248_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_248_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_249_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_249_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_249_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_249_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_250_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_250_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_250_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_250_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_251_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_251_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_251_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_251_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_252_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_252_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_252_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_252_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_253_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_253_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_253_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_253_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_254_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_254_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_254_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_254_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_255_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_255_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_255_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_255_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_256_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_256_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_256_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_256_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_257_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_257_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_257_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_257_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_258_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_258_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_258_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_258_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_259_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_259_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_259_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_259_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_260_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_260_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_260_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_260_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_261_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_261_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_261_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_261_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_262_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_262_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_262_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_262_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_263_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_263_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_263_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_263_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_264_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_264_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_264_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_264_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_265_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_265_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_265_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_265_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_266_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_266_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_266_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_266_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_267_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_267_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_267_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_267_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_268_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_268_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_268_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_268_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_269_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_269_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_269_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_269_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_270_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_270_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_270_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_270_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_271_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_271_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_271_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_271_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_272_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_272_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_272_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_272_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_273_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_273_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_273_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_273_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_274_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_274_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_274_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_274_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_275_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_275_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_275_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_275_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_276_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_276_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_276_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_276_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_277_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_277_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_277_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_277_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_278_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_278_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_278_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_278_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_279_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_279_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_279_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_279_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_280_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_280_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_280_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_280_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_281_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_281_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_281_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_281_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_282_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_282_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_282_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_282_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_283_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_283_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_283_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_283_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_284_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_284_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_284_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_284_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_285_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_285_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_285_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_285_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_286_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_286_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_286_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_286_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_287_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_287_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_287_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_287_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_288_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_288_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_288_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_288_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_289_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_289_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_289_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_289_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_290_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_290_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_290_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_290_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_291_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_291_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_291_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_291_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_292_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_292_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_292_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_292_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_293_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_293_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_293_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_293_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_294_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_294_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_294_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_294_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_295_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_295_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_295_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_295_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_296_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_296_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_296_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_296_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_297_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_297_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_297_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_297_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_298_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_298_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_298_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_298_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_299_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_299_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_299_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_299_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_300_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_300_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_300_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_300_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_301_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_301_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_301_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_301_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_302_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_302_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_302_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_302_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_303_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_303_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_303_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_303_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_304_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_304_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_304_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_304_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_305_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_305_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_305_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_305_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_306_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_306_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_306_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_306_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_307_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_307_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_307_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_307_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_308_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_308_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_308_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_308_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_309_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_309_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_309_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_309_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_310_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_310_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_310_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_310_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_311_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_311_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_311_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_311_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_312_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_312_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_312_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_312_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_313_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_313_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_313_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_313_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_314_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_314_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_314_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_314_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_315_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_315_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_315_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_315_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_316_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_316_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_316_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_316_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_317_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_317_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_317_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_317_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_318_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_318_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_318_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_318_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_319_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_319_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_319_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_319_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_320_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_320_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_320_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_320_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_321_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_321_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_321_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_321_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_322_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_322_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_322_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_322_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_323_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_323_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_323_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_323_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_324_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_324_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_324_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_324_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_325_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_325_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_325_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_325_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_326_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_326_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_326_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_326_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_327_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_327_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_327_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_327_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_328_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_328_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_328_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_328_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_329_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_329_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_329_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_329_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_330_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_330_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_330_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_330_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_331_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_331_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_331_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_331_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_332_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_332_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_332_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_332_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_333_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_333_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_333_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_333_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_334_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_334_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_334_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_334_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_335_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_335_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_335_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_335_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_336_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_336_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_336_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_336_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_337_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_337_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_337_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_337_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_338_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_338_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_338_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_338_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_339_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_339_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_339_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_339_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_340_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_340_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_340_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_340_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_341_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_341_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_341_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_341_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_342_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_342_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_342_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_342_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_343_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_343_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_343_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_343_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_344_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_344_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_344_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_344_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_345_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_345_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_345_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_345_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_346_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_346_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_346_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_346_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_347_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_347_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_347_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_347_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_348_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_348_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_348_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_348_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_349_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_349_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_349_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_349_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_350_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_350_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_350_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_350_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_351_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_351_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_351_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_351_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_352_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_352_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_352_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_352_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_353_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_353_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_353_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_353_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_354_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_354_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_354_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_354_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_355_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_355_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_355_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_355_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_356_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_356_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_356_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_356_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_357_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_357_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_357_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_357_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_358_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_358_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_358_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_358_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_359_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_359_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_359_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_359_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_360_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_360_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_360_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_360_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_361_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_361_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_361_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_361_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_362_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_362_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_362_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_362_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_363_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_363_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_363_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_363_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_364_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_364_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_364_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_364_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_365_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_365_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_365_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_365_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_366_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_366_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_366_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_366_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_367_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_367_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_367_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_367_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_368_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_368_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_368_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_368_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_369_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_369_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_369_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_369_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_370_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_370_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_370_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_370_io_value; // @[coverage.scala 107:33]
  wire  SaturatingCounter_371_clock; // @[coverage.scala 105:33]
  wire  SaturatingCounter_371_reset; // @[coverage.scala 105:33]
  wire  SaturatingCounter_371_io_enable; // @[coverage.scala 105:33]
  wire  SaturatingCounter_371_io_value; // @[coverage.scala 105:33]
  wire  SaturatingCounter_372_clock; // @[coverage.scala 107:33]
  wire  SaturatingCounter_372_reset; // @[coverage.scala 107:33]
  wire  SaturatingCounter_372_io_enable; // @[coverage.scala 107:33]
  wire  SaturatingCounter_372_io_value; // @[coverage.scala 107:33]
  wire [63:0] input_bytes = {io_input_bytes_0,io_input_bytes_1,io_input_bytes_2,io_input_bytes_3,io_input_bytes_4,io_input_bytes_5,io_input_bytes_6,io_input_bytes_7}; // @[Cat.scala 29:58]
  wire [6:0] _T_12 = {6'h0,SaturatingCounter_1_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_16 = {6'h0,SaturatingCounter_3_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_20 = {6'h0,SaturatingCounter_5_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_24 = {6'h0,SaturatingCounter_7_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_28 = {6'h0,SaturatingCounter_9_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_32 = {6'h0,SaturatingCounter_11_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_36 = {6'h0,SaturatingCounter_13_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_40 = {6'h0,SaturatingCounter_15_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_44 = {6'h0,SaturatingCounter_17_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_48 = {6'h0,SaturatingCounter_19_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_52 = {6'h0,SaturatingCounter_21_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_56 = {6'h0,SaturatingCounter_23_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_60 = {6'h0,SaturatingCounter_25_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_64 = {6'h0,SaturatingCounter_27_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_68 = {6'h0,SaturatingCounter_29_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_72 = {6'h0,SaturatingCounter_31_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_76 = {6'h0,SaturatingCounter_33_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_80 = {6'h0,SaturatingCounter_35_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_84 = {6'h0,SaturatingCounter_37_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_88 = {6'h0,SaturatingCounter_39_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_92 = {6'h0,SaturatingCounter_41_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_96 = {6'h0,SaturatingCounter_43_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_100 = {6'h0,SaturatingCounter_45_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_104 = {6'h0,SaturatingCounter_47_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_108 = {6'h0,SaturatingCounter_49_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_112 = {6'h0,SaturatingCounter_51_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_116 = {6'h0,SaturatingCounter_53_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_120 = {6'h0,SaturatingCounter_55_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_124 = {6'h0,SaturatingCounter_57_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_128 = {6'h0,SaturatingCounter_59_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_132 = {6'h0,SaturatingCounter_61_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_136 = {6'h0,SaturatingCounter_63_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_140 = {6'h0,SaturatingCounter_65_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_144 = {6'h0,SaturatingCounter_67_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_148 = {6'h0,SaturatingCounter_69_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_152 = {6'h0,SaturatingCounter_71_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_156 = {6'h0,SaturatingCounter_73_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_160 = {6'h0,SaturatingCounter_75_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_164 = {6'h0,SaturatingCounter_77_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_168 = {6'h0,SaturatingCounter_79_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_172 = {6'h0,SaturatingCounter_81_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_176 = {6'h0,SaturatingCounter_83_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_180 = {6'h0,SaturatingCounter_85_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_184 = {6'h0,SaturatingCounter_87_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_188 = {6'h0,SaturatingCounter_89_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_192 = {6'h0,SaturatingCounter_91_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_196 = {6'h0,SaturatingCounter_93_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_200 = {6'h0,SaturatingCounter_95_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_204 = {6'h0,SaturatingCounter_97_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_208 = {6'h0,SaturatingCounter_99_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_212 = {6'h0,SaturatingCounter_101_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_216 = {6'h0,SaturatingCounter_103_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_220 = {6'h0,SaturatingCounter_105_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_224 = {6'h0,SaturatingCounter_107_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_228 = {6'h0,SaturatingCounter_109_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_232 = {6'h0,SaturatingCounter_111_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_236 = {6'h0,SaturatingCounter_113_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_240 = {6'h0,SaturatingCounter_115_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_244 = {6'h0,SaturatingCounter_117_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_248 = {6'h0,SaturatingCounter_119_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_252 = {6'h0,SaturatingCounter_121_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_256 = {6'h0,SaturatingCounter_123_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_260 = {6'h0,SaturatingCounter_125_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_264 = {6'h0,SaturatingCounter_127_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_268 = {6'h0,SaturatingCounter_129_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_272 = {6'h0,SaturatingCounter_131_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_276 = {6'h0,SaturatingCounter_133_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_280 = {6'h0,SaturatingCounter_135_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_284 = {6'h0,SaturatingCounter_137_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_288 = {6'h0,SaturatingCounter_139_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_292 = {6'h0,SaturatingCounter_141_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_296 = {6'h0,SaturatingCounter_143_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_300 = {6'h0,SaturatingCounter_145_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_304 = {6'h0,SaturatingCounter_147_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_308 = {6'h0,SaturatingCounter_149_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_312 = {6'h0,SaturatingCounter_151_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_316 = {6'h0,SaturatingCounter_153_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_320 = {6'h0,SaturatingCounter_155_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_324 = {6'h0,SaturatingCounter_157_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_328 = {6'h0,SaturatingCounter_159_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_332 = {6'h0,SaturatingCounter_161_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_336 = {6'h0,SaturatingCounter_163_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_340 = {6'h0,SaturatingCounter_165_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_344 = {6'h0,SaturatingCounter_167_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_348 = {6'h0,SaturatingCounter_169_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_352 = {6'h0,SaturatingCounter_171_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_356 = {6'h0,SaturatingCounter_173_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_360 = {6'h0,SaturatingCounter_175_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_364 = {6'h0,SaturatingCounter_177_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_368 = {6'h0,SaturatingCounter_179_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_372 = {6'h0,SaturatingCounter_181_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_376 = {6'h0,SaturatingCounter_183_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_380 = {6'h0,SaturatingCounter_185_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_384 = {6'h0,SaturatingCounter_187_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_388 = {6'h0,SaturatingCounter_189_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_392 = {6'h0,SaturatingCounter_191_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_396 = {6'h0,SaturatingCounter_193_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_400 = {6'h0,SaturatingCounter_195_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_404 = {6'h0,SaturatingCounter_197_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_408 = {6'h0,SaturatingCounter_199_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_412 = {6'h0,SaturatingCounter_201_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_416 = {6'h0,SaturatingCounter_203_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_420 = {6'h0,SaturatingCounter_205_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_424 = {6'h0,SaturatingCounter_207_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_428 = {6'h0,SaturatingCounter_209_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_432 = {6'h0,SaturatingCounter_211_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_436 = {6'h0,SaturatingCounter_213_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_440 = {6'h0,SaturatingCounter_215_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_444 = {6'h0,SaturatingCounter_217_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_448 = {6'h0,SaturatingCounter_219_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_452 = {6'h0,SaturatingCounter_221_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_456 = {6'h0,SaturatingCounter_223_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_460 = {6'h0,SaturatingCounter_225_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_464 = {6'h0,SaturatingCounter_227_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_468 = {6'h0,SaturatingCounter_229_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_472 = {6'h0,SaturatingCounter_231_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_476 = {6'h0,SaturatingCounter_233_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_480 = {6'h0,SaturatingCounter_235_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_484 = {6'h0,SaturatingCounter_237_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_488 = {6'h0,SaturatingCounter_239_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_492 = {6'h0,SaturatingCounter_241_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_496 = {6'h0,SaturatingCounter_243_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_500 = {6'h0,SaturatingCounter_245_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_504 = {6'h0,SaturatingCounter_247_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_508 = {6'h0,SaturatingCounter_249_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_512 = {6'h0,SaturatingCounter_251_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_516 = {6'h0,SaturatingCounter_253_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_520 = {6'h0,SaturatingCounter_255_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_524 = {6'h0,SaturatingCounter_257_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_528 = {6'h0,SaturatingCounter_259_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_532 = {6'h0,SaturatingCounter_261_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_536 = {6'h0,SaturatingCounter_263_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_540 = {6'h0,SaturatingCounter_265_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_544 = {6'h0,SaturatingCounter_267_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_548 = {6'h0,SaturatingCounter_269_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_552 = {6'h0,SaturatingCounter_271_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_556 = {6'h0,SaturatingCounter_273_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_560 = {6'h0,SaturatingCounter_275_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_564 = {6'h0,SaturatingCounter_277_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_568 = {6'h0,SaturatingCounter_279_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_572 = {6'h0,SaturatingCounter_281_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_576 = {6'h0,SaturatingCounter_283_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_580 = {6'h0,SaturatingCounter_285_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_584 = {6'h0,SaturatingCounter_287_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_588 = {6'h0,SaturatingCounter_289_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_592 = {6'h0,SaturatingCounter_291_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_596 = {6'h0,SaturatingCounter_293_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_600 = {6'h0,SaturatingCounter_295_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_604 = {6'h0,SaturatingCounter_297_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_608 = {6'h0,SaturatingCounter_299_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_612 = {6'h0,SaturatingCounter_301_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_616 = {6'h0,SaturatingCounter_303_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_620 = {6'h0,SaturatingCounter_305_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_624 = {6'h0,SaturatingCounter_307_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_628 = {6'h0,SaturatingCounter_309_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_632 = {6'h0,SaturatingCounter_311_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_636 = {6'h0,SaturatingCounter_313_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_640 = {6'h0,SaturatingCounter_315_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_644 = {6'h0,SaturatingCounter_317_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_648 = {6'h0,SaturatingCounter_319_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_652 = {6'h0,SaturatingCounter_321_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_656 = {6'h0,SaturatingCounter_323_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_660 = {6'h0,SaturatingCounter_325_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_664 = {6'h0,SaturatingCounter_327_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_668 = {6'h0,SaturatingCounter_329_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_672 = {6'h0,SaturatingCounter_331_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_676 = {6'h0,SaturatingCounter_333_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_680 = {6'h0,SaturatingCounter_335_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_684 = {6'h0,SaturatingCounter_337_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_688 = {6'h0,SaturatingCounter_339_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_692 = {6'h0,SaturatingCounter_341_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_696 = {6'h0,SaturatingCounter_343_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_700 = {6'h0,SaturatingCounter_345_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_704 = {6'h0,SaturatingCounter_347_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_708 = {6'h0,SaturatingCounter_349_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_712 = {6'h0,SaturatingCounter_351_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_716 = {6'h0,SaturatingCounter_353_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_720 = {6'h0,SaturatingCounter_355_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_724 = {6'h0,SaturatingCounter_357_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_728 = {6'h0,SaturatingCounter_359_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_732 = {6'h0,SaturatingCounter_361_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_736 = {6'h0,SaturatingCounter_363_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_740 = {6'h0,SaturatingCounter_365_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_744 = {6'h0,SaturatingCounter_367_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_748 = {6'h0,SaturatingCounter_369_io_value}; // @[Cat.scala 29:58]
  wire [6:0] _T_752 = {6'h0,SaturatingCounter_371_io_value}; // @[Cat.scala 29:58]
  DUT dut ( // @[VerilatorHarness.scala 42:25]
    .clock(dut_clock),
    .reset(dut_reset),
    .io_meta_reset(dut_io_meta_reset),
    .io_inputs(dut_io_inputs),
    .io_coverage_0(dut_io_coverage_0),
    .io_coverage_1(dut_io_coverage_1),
    .io_coverage_2(dut_io_coverage_2),
    .io_coverage_3(dut_io_coverage_3),
    .io_coverage_4(dut_io_coverage_4),
    .io_coverage_5(dut_io_coverage_5),
    .io_coverage_6(dut_io_coverage_6),
    .io_coverage_7(dut_io_coverage_7),
    .io_coverage_8(dut_io_coverage_8),
    .io_coverage_9(dut_io_coverage_9),
    .io_coverage_10(dut_io_coverage_10),
    .io_coverage_11(dut_io_coverage_11),
    .io_coverage_12(dut_io_coverage_12),
    .io_coverage_13(dut_io_coverage_13),
    .io_coverage_14(dut_io_coverage_14),
    .io_coverage_15(dut_io_coverage_15),
    .io_coverage_16(dut_io_coverage_16),
    .io_coverage_17(dut_io_coverage_17),
    .io_coverage_18(dut_io_coverage_18),
    .io_coverage_19(dut_io_coverage_19),
    .io_coverage_20(dut_io_coverage_20),
    .io_coverage_21(dut_io_coverage_21),
    .io_coverage_22(dut_io_coverage_22),
    .io_coverage_23(dut_io_coverage_23),
    .io_coverage_24(dut_io_coverage_24),
    .io_coverage_25(dut_io_coverage_25),
    .io_coverage_26(dut_io_coverage_26),
    .io_coverage_27(dut_io_coverage_27),
    .io_coverage_28(dut_io_coverage_28),
    .io_coverage_29(dut_io_coverage_29),
    .io_coverage_30(dut_io_coverage_30),
    .io_coverage_31(dut_io_coverage_31),
    .io_coverage_32(dut_io_coverage_32),
    .io_coverage_33(dut_io_coverage_33),
    .io_coverage_34(dut_io_coverage_34),
    .io_coverage_35(dut_io_coverage_35),
    .io_coverage_36(dut_io_coverage_36),
    .io_coverage_37(dut_io_coverage_37),
    .io_coverage_38(dut_io_coverage_38),
    .io_coverage_39(dut_io_coverage_39),
    .io_coverage_40(dut_io_coverage_40),
    .io_coverage_41(dut_io_coverage_41),
    .io_coverage_42(dut_io_coverage_42),
    .io_coverage_43(dut_io_coverage_43),
    .io_coverage_44(dut_io_coverage_44),
    .io_coverage_45(dut_io_coverage_45),
    .io_coverage_46(dut_io_coverage_46),
    .io_coverage_47(dut_io_coverage_47),
    .io_coverage_48(dut_io_coverage_48),
    .io_coverage_49(dut_io_coverage_49),
    .io_coverage_50(dut_io_coverage_50),
    .io_coverage_51(dut_io_coverage_51),
    .io_coverage_52(dut_io_coverage_52),
    .io_coverage_53(dut_io_coverage_53),
    .io_coverage_54(dut_io_coverage_54),
    .io_coverage_55(dut_io_coverage_55),
    .io_coverage_56(dut_io_coverage_56),
    .io_coverage_57(dut_io_coverage_57),
    .io_coverage_58(dut_io_coverage_58),
    .io_coverage_59(dut_io_coverage_59),
    .io_coverage_60(dut_io_coverage_60),
    .io_coverage_61(dut_io_coverage_61),
    .io_coverage_62(dut_io_coverage_62),
    .io_coverage_63(dut_io_coverage_63),
    .io_coverage_64(dut_io_coverage_64),
    .io_coverage_65(dut_io_coverage_65),
    .io_coverage_66(dut_io_coverage_66),
    .io_coverage_67(dut_io_coverage_67),
    .io_coverage_68(dut_io_coverage_68),
    .io_coverage_69(dut_io_coverage_69),
    .io_coverage_70(dut_io_coverage_70),
    .io_coverage_71(dut_io_coverage_71),
    .io_coverage_72(dut_io_coverage_72),
    .io_coverage_73(dut_io_coverage_73),
    .io_coverage_74(dut_io_coverage_74),
    .io_coverage_75(dut_io_coverage_75),
    .io_coverage_76(dut_io_coverage_76),
    .io_coverage_77(dut_io_coverage_77),
    .io_coverage_78(dut_io_coverage_78),
    .io_coverage_79(dut_io_coverage_79),
    .io_coverage_80(dut_io_coverage_80),
    .io_coverage_81(dut_io_coverage_81),
    .io_coverage_82(dut_io_coverage_82),
    .io_coverage_83(dut_io_coverage_83),
    .io_coverage_84(dut_io_coverage_84),
    .io_coverage_85(dut_io_coverage_85),
    .io_coverage_86(dut_io_coverage_86),
    .io_coverage_87(dut_io_coverage_87),
    .io_coverage_88(dut_io_coverage_88),
    .io_coverage_89(dut_io_coverage_89),
    .io_coverage_90(dut_io_coverage_90),
    .io_coverage_91(dut_io_coverage_91),
    .io_coverage_92(dut_io_coverage_92),
    .io_coverage_93(dut_io_coverage_93),
    .io_coverage_94(dut_io_coverage_94),
    .io_coverage_95(dut_io_coverage_95),
    .io_coverage_96(dut_io_coverage_96),
    .io_coverage_97(dut_io_coverage_97),
    .io_coverage_98(dut_io_coverage_98),
    .io_coverage_99(dut_io_coverage_99),
    .io_coverage_100(dut_io_coverage_100),
    .io_coverage_101(dut_io_coverage_101),
    .io_coverage_102(dut_io_coverage_102),
    .io_coverage_103(dut_io_coverage_103),
    .io_coverage_104(dut_io_coverage_104),
    .io_coverage_105(dut_io_coverage_105),
    .io_coverage_106(dut_io_coverage_106),
    .io_coverage_107(dut_io_coverage_107),
    .io_coverage_108(dut_io_coverage_108),
    .io_coverage_109(dut_io_coverage_109),
    .io_coverage_110(dut_io_coverage_110),
    .io_coverage_111(dut_io_coverage_111),
    .io_coverage_112(dut_io_coverage_112),
    .io_coverage_113(dut_io_coverage_113),
    .io_coverage_114(dut_io_coverage_114),
    .io_coverage_115(dut_io_coverage_115),
    .io_coverage_116(dut_io_coverage_116),
    .io_coverage_117(dut_io_coverage_117),
    .io_coverage_118(dut_io_coverage_118),
    .io_coverage_119(dut_io_coverage_119),
    .io_coverage_120(dut_io_coverage_120),
    .io_coverage_121(dut_io_coverage_121),
    .io_coverage_122(dut_io_coverage_122),
    .io_coverage_123(dut_io_coverage_123),
    .io_coverage_124(dut_io_coverage_124),
    .io_coverage_125(dut_io_coverage_125),
    .io_coverage_126(dut_io_coverage_126),
    .io_coverage_127(dut_io_coverage_127),
    .io_coverage_128(dut_io_coverage_128),
    .io_coverage_129(dut_io_coverage_129),
    .io_coverage_130(dut_io_coverage_130),
    .io_coverage_131(dut_io_coverage_131),
    .io_coverage_132(dut_io_coverage_132),
    .io_coverage_133(dut_io_coverage_133),
    .io_coverage_134(dut_io_coverage_134),
    .io_coverage_135(dut_io_coverage_135),
    .io_coverage_136(dut_io_coverage_136),
    .io_coverage_137(dut_io_coverage_137),
    .io_coverage_138(dut_io_coverage_138),
    .io_coverage_139(dut_io_coverage_139),
    .io_coverage_140(dut_io_coverage_140),
    .io_coverage_141(dut_io_coverage_141),
    .io_coverage_142(dut_io_coverage_142),
    .io_coverage_143(dut_io_coverage_143),
    .io_coverage_144(dut_io_coverage_144),
    .io_coverage_145(dut_io_coverage_145),
    .io_coverage_146(dut_io_coverage_146),
    .io_coverage_147(dut_io_coverage_147),
    .io_coverage_148(dut_io_coverage_148),
    .io_coverage_149(dut_io_coverage_149),
    .io_coverage_150(dut_io_coverage_150),
    .io_coverage_151(dut_io_coverage_151),
    .io_coverage_152(dut_io_coverage_152),
    .io_coverage_153(dut_io_coverage_153),
    .io_coverage_154(dut_io_coverage_154),
    .io_coverage_155(dut_io_coverage_155),
    .io_coverage_156(dut_io_coverage_156),
    .io_coverage_157(dut_io_coverage_157),
    .io_coverage_158(dut_io_coverage_158),
    .io_coverage_159(dut_io_coverage_159),
    .io_coverage_160(dut_io_coverage_160),
    .io_coverage_161(dut_io_coverage_161),
    .io_coverage_162(dut_io_coverage_162),
    .io_coverage_163(dut_io_coverage_163),
    .io_coverage_164(dut_io_coverage_164),
    .io_coverage_165(dut_io_coverage_165),
    .io_coverage_166(dut_io_coverage_166),
    .io_coverage_167(dut_io_coverage_167),
    .io_coverage_168(dut_io_coverage_168),
    .io_coverage_169(dut_io_coverage_169),
    .io_coverage_170(dut_io_coverage_170),
    .io_coverage_171(dut_io_coverage_171),
    .io_coverage_172(dut_io_coverage_172),
    .io_coverage_173(dut_io_coverage_173),
    .io_coverage_174(dut_io_coverage_174),
    .io_coverage_175(dut_io_coverage_175),
    .io_coverage_176(dut_io_coverage_176),
    .io_coverage_177(dut_io_coverage_177),
    .io_coverage_178(dut_io_coverage_178),
    .io_coverage_179(dut_io_coverage_179),
    .io_coverage_180(dut_io_coverage_180),
    .io_coverage_181(dut_io_coverage_181),
    .io_coverage_182(dut_io_coverage_182),
    .io_coverage_183(dut_io_coverage_183),
    .io_coverage_184(dut_io_coverage_184),
    .io_coverage_185(dut_io_coverage_185),
    .io_coverage_186(dut_io_coverage_186)
  );
  SaturatingCounter SaturatingCounter ( // @[coverage.scala 121:35]
    .clock(SaturatingCounter_clock),
    .reset(SaturatingCounter_reset),
    .io_enable(SaturatingCounter_io_enable),
    .io_value(SaturatingCounter_io_value)
  );
  SaturatingCounter SaturatingCounter_1 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_1_clock),
    .reset(SaturatingCounter_1_reset),
    .io_enable(SaturatingCounter_1_io_enable),
    .io_value(SaturatingCounter_1_io_value)
  );
  SaturatingCounter SaturatingCounter_2 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_2_clock),
    .reset(SaturatingCounter_2_reset),
    .io_enable(SaturatingCounter_2_io_enable),
    .io_value(SaturatingCounter_2_io_value)
  );
  SaturatingCounter SaturatingCounter_3 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_3_clock),
    .reset(SaturatingCounter_3_reset),
    .io_enable(SaturatingCounter_3_io_enable),
    .io_value(SaturatingCounter_3_io_value)
  );
  SaturatingCounter SaturatingCounter_4 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_4_clock),
    .reset(SaturatingCounter_4_reset),
    .io_enable(SaturatingCounter_4_io_enable),
    .io_value(SaturatingCounter_4_io_value)
  );
  SaturatingCounter SaturatingCounter_5 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_5_clock),
    .reset(SaturatingCounter_5_reset),
    .io_enable(SaturatingCounter_5_io_enable),
    .io_value(SaturatingCounter_5_io_value)
  );
  SaturatingCounter SaturatingCounter_6 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_6_clock),
    .reset(SaturatingCounter_6_reset),
    .io_enable(SaturatingCounter_6_io_enable),
    .io_value(SaturatingCounter_6_io_value)
  );
  SaturatingCounter SaturatingCounter_7 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_7_clock),
    .reset(SaturatingCounter_7_reset),
    .io_enable(SaturatingCounter_7_io_enable),
    .io_value(SaturatingCounter_7_io_value)
  );
  SaturatingCounter SaturatingCounter_8 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_8_clock),
    .reset(SaturatingCounter_8_reset),
    .io_enable(SaturatingCounter_8_io_enable),
    .io_value(SaturatingCounter_8_io_value)
  );
  SaturatingCounter SaturatingCounter_9 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_9_clock),
    .reset(SaturatingCounter_9_reset),
    .io_enable(SaturatingCounter_9_io_enable),
    .io_value(SaturatingCounter_9_io_value)
  );
  SaturatingCounter SaturatingCounter_10 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_10_clock),
    .reset(SaturatingCounter_10_reset),
    .io_enable(SaturatingCounter_10_io_enable),
    .io_value(SaturatingCounter_10_io_value)
  );
  SaturatingCounter SaturatingCounter_11 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_11_clock),
    .reset(SaturatingCounter_11_reset),
    .io_enable(SaturatingCounter_11_io_enable),
    .io_value(SaturatingCounter_11_io_value)
  );
  SaturatingCounter SaturatingCounter_12 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_12_clock),
    .reset(SaturatingCounter_12_reset),
    .io_enable(SaturatingCounter_12_io_enable),
    .io_value(SaturatingCounter_12_io_value)
  );
  SaturatingCounter SaturatingCounter_13 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_13_clock),
    .reset(SaturatingCounter_13_reset),
    .io_enable(SaturatingCounter_13_io_enable),
    .io_value(SaturatingCounter_13_io_value)
  );
  SaturatingCounter SaturatingCounter_14 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_14_clock),
    .reset(SaturatingCounter_14_reset),
    .io_enable(SaturatingCounter_14_io_enable),
    .io_value(SaturatingCounter_14_io_value)
  );
  SaturatingCounter SaturatingCounter_15 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_15_clock),
    .reset(SaturatingCounter_15_reset),
    .io_enable(SaturatingCounter_15_io_enable),
    .io_value(SaturatingCounter_15_io_value)
  );
  SaturatingCounter SaturatingCounter_16 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_16_clock),
    .reset(SaturatingCounter_16_reset),
    .io_enable(SaturatingCounter_16_io_enable),
    .io_value(SaturatingCounter_16_io_value)
  );
  SaturatingCounter SaturatingCounter_17 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_17_clock),
    .reset(SaturatingCounter_17_reset),
    .io_enable(SaturatingCounter_17_io_enable),
    .io_value(SaturatingCounter_17_io_value)
  );
  SaturatingCounter SaturatingCounter_18 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_18_clock),
    .reset(SaturatingCounter_18_reset),
    .io_enable(SaturatingCounter_18_io_enable),
    .io_value(SaturatingCounter_18_io_value)
  );
  SaturatingCounter SaturatingCounter_19 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_19_clock),
    .reset(SaturatingCounter_19_reset),
    .io_enable(SaturatingCounter_19_io_enable),
    .io_value(SaturatingCounter_19_io_value)
  );
  SaturatingCounter SaturatingCounter_20 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_20_clock),
    .reset(SaturatingCounter_20_reset),
    .io_enable(SaturatingCounter_20_io_enable),
    .io_value(SaturatingCounter_20_io_value)
  );
  SaturatingCounter SaturatingCounter_21 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_21_clock),
    .reset(SaturatingCounter_21_reset),
    .io_enable(SaturatingCounter_21_io_enable),
    .io_value(SaturatingCounter_21_io_value)
  );
  SaturatingCounter SaturatingCounter_22 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_22_clock),
    .reset(SaturatingCounter_22_reset),
    .io_enable(SaturatingCounter_22_io_enable),
    .io_value(SaturatingCounter_22_io_value)
  );
  SaturatingCounter SaturatingCounter_23 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_23_clock),
    .reset(SaturatingCounter_23_reset),
    .io_enable(SaturatingCounter_23_io_enable),
    .io_value(SaturatingCounter_23_io_value)
  );
  SaturatingCounter SaturatingCounter_24 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_24_clock),
    .reset(SaturatingCounter_24_reset),
    .io_enable(SaturatingCounter_24_io_enable),
    .io_value(SaturatingCounter_24_io_value)
  );
  SaturatingCounter SaturatingCounter_25 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_25_clock),
    .reset(SaturatingCounter_25_reset),
    .io_enable(SaturatingCounter_25_io_enable),
    .io_value(SaturatingCounter_25_io_value)
  );
  SaturatingCounter SaturatingCounter_26 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_26_clock),
    .reset(SaturatingCounter_26_reset),
    .io_enable(SaturatingCounter_26_io_enable),
    .io_value(SaturatingCounter_26_io_value)
  );
  SaturatingCounter SaturatingCounter_27 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_27_clock),
    .reset(SaturatingCounter_27_reset),
    .io_enable(SaturatingCounter_27_io_enable),
    .io_value(SaturatingCounter_27_io_value)
  );
  SaturatingCounter SaturatingCounter_28 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_28_clock),
    .reset(SaturatingCounter_28_reset),
    .io_enable(SaturatingCounter_28_io_enable),
    .io_value(SaturatingCounter_28_io_value)
  );
  SaturatingCounter SaturatingCounter_29 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_29_clock),
    .reset(SaturatingCounter_29_reset),
    .io_enable(SaturatingCounter_29_io_enable),
    .io_value(SaturatingCounter_29_io_value)
  );
  SaturatingCounter SaturatingCounter_30 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_30_clock),
    .reset(SaturatingCounter_30_reset),
    .io_enable(SaturatingCounter_30_io_enable),
    .io_value(SaturatingCounter_30_io_value)
  );
  SaturatingCounter SaturatingCounter_31 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_31_clock),
    .reset(SaturatingCounter_31_reset),
    .io_enable(SaturatingCounter_31_io_enable),
    .io_value(SaturatingCounter_31_io_value)
  );
  SaturatingCounter SaturatingCounter_32 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_32_clock),
    .reset(SaturatingCounter_32_reset),
    .io_enable(SaturatingCounter_32_io_enable),
    .io_value(SaturatingCounter_32_io_value)
  );
  SaturatingCounter SaturatingCounter_33 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_33_clock),
    .reset(SaturatingCounter_33_reset),
    .io_enable(SaturatingCounter_33_io_enable),
    .io_value(SaturatingCounter_33_io_value)
  );
  SaturatingCounter SaturatingCounter_34 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_34_clock),
    .reset(SaturatingCounter_34_reset),
    .io_enable(SaturatingCounter_34_io_enable),
    .io_value(SaturatingCounter_34_io_value)
  );
  SaturatingCounter SaturatingCounter_35 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_35_clock),
    .reset(SaturatingCounter_35_reset),
    .io_enable(SaturatingCounter_35_io_enable),
    .io_value(SaturatingCounter_35_io_value)
  );
  SaturatingCounter SaturatingCounter_36 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_36_clock),
    .reset(SaturatingCounter_36_reset),
    .io_enable(SaturatingCounter_36_io_enable),
    .io_value(SaturatingCounter_36_io_value)
  );
  SaturatingCounter SaturatingCounter_37 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_37_clock),
    .reset(SaturatingCounter_37_reset),
    .io_enable(SaturatingCounter_37_io_enable),
    .io_value(SaturatingCounter_37_io_value)
  );
  SaturatingCounter SaturatingCounter_38 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_38_clock),
    .reset(SaturatingCounter_38_reset),
    .io_enable(SaturatingCounter_38_io_enable),
    .io_value(SaturatingCounter_38_io_value)
  );
  SaturatingCounter SaturatingCounter_39 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_39_clock),
    .reset(SaturatingCounter_39_reset),
    .io_enable(SaturatingCounter_39_io_enable),
    .io_value(SaturatingCounter_39_io_value)
  );
  SaturatingCounter SaturatingCounter_40 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_40_clock),
    .reset(SaturatingCounter_40_reset),
    .io_enable(SaturatingCounter_40_io_enable),
    .io_value(SaturatingCounter_40_io_value)
  );
  SaturatingCounter SaturatingCounter_41 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_41_clock),
    .reset(SaturatingCounter_41_reset),
    .io_enable(SaturatingCounter_41_io_enable),
    .io_value(SaturatingCounter_41_io_value)
  );
  SaturatingCounter SaturatingCounter_42 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_42_clock),
    .reset(SaturatingCounter_42_reset),
    .io_enable(SaturatingCounter_42_io_enable),
    .io_value(SaturatingCounter_42_io_value)
  );
  SaturatingCounter SaturatingCounter_43 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_43_clock),
    .reset(SaturatingCounter_43_reset),
    .io_enable(SaturatingCounter_43_io_enable),
    .io_value(SaturatingCounter_43_io_value)
  );
  SaturatingCounter SaturatingCounter_44 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_44_clock),
    .reset(SaturatingCounter_44_reset),
    .io_enable(SaturatingCounter_44_io_enable),
    .io_value(SaturatingCounter_44_io_value)
  );
  SaturatingCounter SaturatingCounter_45 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_45_clock),
    .reset(SaturatingCounter_45_reset),
    .io_enable(SaturatingCounter_45_io_enable),
    .io_value(SaturatingCounter_45_io_value)
  );
  SaturatingCounter SaturatingCounter_46 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_46_clock),
    .reset(SaturatingCounter_46_reset),
    .io_enable(SaturatingCounter_46_io_enable),
    .io_value(SaturatingCounter_46_io_value)
  );
  SaturatingCounter SaturatingCounter_47 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_47_clock),
    .reset(SaturatingCounter_47_reset),
    .io_enable(SaturatingCounter_47_io_enable),
    .io_value(SaturatingCounter_47_io_value)
  );
  SaturatingCounter SaturatingCounter_48 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_48_clock),
    .reset(SaturatingCounter_48_reset),
    .io_enable(SaturatingCounter_48_io_enable),
    .io_value(SaturatingCounter_48_io_value)
  );
  SaturatingCounter SaturatingCounter_49 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_49_clock),
    .reset(SaturatingCounter_49_reset),
    .io_enable(SaturatingCounter_49_io_enable),
    .io_value(SaturatingCounter_49_io_value)
  );
  SaturatingCounter SaturatingCounter_50 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_50_clock),
    .reset(SaturatingCounter_50_reset),
    .io_enable(SaturatingCounter_50_io_enable),
    .io_value(SaturatingCounter_50_io_value)
  );
  SaturatingCounter SaturatingCounter_51 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_51_clock),
    .reset(SaturatingCounter_51_reset),
    .io_enable(SaturatingCounter_51_io_enable),
    .io_value(SaturatingCounter_51_io_value)
  );
  SaturatingCounter SaturatingCounter_52 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_52_clock),
    .reset(SaturatingCounter_52_reset),
    .io_enable(SaturatingCounter_52_io_enable),
    .io_value(SaturatingCounter_52_io_value)
  );
  SaturatingCounter SaturatingCounter_53 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_53_clock),
    .reset(SaturatingCounter_53_reset),
    .io_enable(SaturatingCounter_53_io_enable),
    .io_value(SaturatingCounter_53_io_value)
  );
  SaturatingCounter SaturatingCounter_54 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_54_clock),
    .reset(SaturatingCounter_54_reset),
    .io_enable(SaturatingCounter_54_io_enable),
    .io_value(SaturatingCounter_54_io_value)
  );
  SaturatingCounter SaturatingCounter_55 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_55_clock),
    .reset(SaturatingCounter_55_reset),
    .io_enable(SaturatingCounter_55_io_enable),
    .io_value(SaturatingCounter_55_io_value)
  );
  SaturatingCounter SaturatingCounter_56 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_56_clock),
    .reset(SaturatingCounter_56_reset),
    .io_enable(SaturatingCounter_56_io_enable),
    .io_value(SaturatingCounter_56_io_value)
  );
  SaturatingCounter SaturatingCounter_57 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_57_clock),
    .reset(SaturatingCounter_57_reset),
    .io_enable(SaturatingCounter_57_io_enable),
    .io_value(SaturatingCounter_57_io_value)
  );
  SaturatingCounter SaturatingCounter_58 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_58_clock),
    .reset(SaturatingCounter_58_reset),
    .io_enable(SaturatingCounter_58_io_enable),
    .io_value(SaturatingCounter_58_io_value)
  );
  SaturatingCounter SaturatingCounter_59 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_59_clock),
    .reset(SaturatingCounter_59_reset),
    .io_enable(SaturatingCounter_59_io_enable),
    .io_value(SaturatingCounter_59_io_value)
  );
  SaturatingCounter SaturatingCounter_60 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_60_clock),
    .reset(SaturatingCounter_60_reset),
    .io_enable(SaturatingCounter_60_io_enable),
    .io_value(SaturatingCounter_60_io_value)
  );
  SaturatingCounter SaturatingCounter_61 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_61_clock),
    .reset(SaturatingCounter_61_reset),
    .io_enable(SaturatingCounter_61_io_enable),
    .io_value(SaturatingCounter_61_io_value)
  );
  SaturatingCounter SaturatingCounter_62 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_62_clock),
    .reset(SaturatingCounter_62_reset),
    .io_enable(SaturatingCounter_62_io_enable),
    .io_value(SaturatingCounter_62_io_value)
  );
  SaturatingCounter SaturatingCounter_63 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_63_clock),
    .reset(SaturatingCounter_63_reset),
    .io_enable(SaturatingCounter_63_io_enable),
    .io_value(SaturatingCounter_63_io_value)
  );
  SaturatingCounter SaturatingCounter_64 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_64_clock),
    .reset(SaturatingCounter_64_reset),
    .io_enable(SaturatingCounter_64_io_enable),
    .io_value(SaturatingCounter_64_io_value)
  );
  SaturatingCounter SaturatingCounter_65 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_65_clock),
    .reset(SaturatingCounter_65_reset),
    .io_enable(SaturatingCounter_65_io_enable),
    .io_value(SaturatingCounter_65_io_value)
  );
  SaturatingCounter SaturatingCounter_66 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_66_clock),
    .reset(SaturatingCounter_66_reset),
    .io_enable(SaturatingCounter_66_io_enable),
    .io_value(SaturatingCounter_66_io_value)
  );
  SaturatingCounter SaturatingCounter_67 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_67_clock),
    .reset(SaturatingCounter_67_reset),
    .io_enable(SaturatingCounter_67_io_enable),
    .io_value(SaturatingCounter_67_io_value)
  );
  SaturatingCounter SaturatingCounter_68 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_68_clock),
    .reset(SaturatingCounter_68_reset),
    .io_enable(SaturatingCounter_68_io_enable),
    .io_value(SaturatingCounter_68_io_value)
  );
  SaturatingCounter SaturatingCounter_69 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_69_clock),
    .reset(SaturatingCounter_69_reset),
    .io_enable(SaturatingCounter_69_io_enable),
    .io_value(SaturatingCounter_69_io_value)
  );
  SaturatingCounter SaturatingCounter_70 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_70_clock),
    .reset(SaturatingCounter_70_reset),
    .io_enable(SaturatingCounter_70_io_enable),
    .io_value(SaturatingCounter_70_io_value)
  );
  SaturatingCounter SaturatingCounter_71 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_71_clock),
    .reset(SaturatingCounter_71_reset),
    .io_enable(SaturatingCounter_71_io_enable),
    .io_value(SaturatingCounter_71_io_value)
  );
  SaturatingCounter SaturatingCounter_72 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_72_clock),
    .reset(SaturatingCounter_72_reset),
    .io_enable(SaturatingCounter_72_io_enable),
    .io_value(SaturatingCounter_72_io_value)
  );
  SaturatingCounter SaturatingCounter_73 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_73_clock),
    .reset(SaturatingCounter_73_reset),
    .io_enable(SaturatingCounter_73_io_enable),
    .io_value(SaturatingCounter_73_io_value)
  );
  SaturatingCounter SaturatingCounter_74 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_74_clock),
    .reset(SaturatingCounter_74_reset),
    .io_enable(SaturatingCounter_74_io_enable),
    .io_value(SaturatingCounter_74_io_value)
  );
  SaturatingCounter SaturatingCounter_75 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_75_clock),
    .reset(SaturatingCounter_75_reset),
    .io_enable(SaturatingCounter_75_io_enable),
    .io_value(SaturatingCounter_75_io_value)
  );
  SaturatingCounter SaturatingCounter_76 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_76_clock),
    .reset(SaturatingCounter_76_reset),
    .io_enable(SaturatingCounter_76_io_enable),
    .io_value(SaturatingCounter_76_io_value)
  );
  SaturatingCounter SaturatingCounter_77 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_77_clock),
    .reset(SaturatingCounter_77_reset),
    .io_enable(SaturatingCounter_77_io_enable),
    .io_value(SaturatingCounter_77_io_value)
  );
  SaturatingCounter SaturatingCounter_78 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_78_clock),
    .reset(SaturatingCounter_78_reset),
    .io_enable(SaturatingCounter_78_io_enable),
    .io_value(SaturatingCounter_78_io_value)
  );
  SaturatingCounter SaturatingCounter_79 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_79_clock),
    .reset(SaturatingCounter_79_reset),
    .io_enable(SaturatingCounter_79_io_enable),
    .io_value(SaturatingCounter_79_io_value)
  );
  SaturatingCounter SaturatingCounter_80 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_80_clock),
    .reset(SaturatingCounter_80_reset),
    .io_enable(SaturatingCounter_80_io_enable),
    .io_value(SaturatingCounter_80_io_value)
  );
  SaturatingCounter SaturatingCounter_81 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_81_clock),
    .reset(SaturatingCounter_81_reset),
    .io_enable(SaturatingCounter_81_io_enable),
    .io_value(SaturatingCounter_81_io_value)
  );
  SaturatingCounter SaturatingCounter_82 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_82_clock),
    .reset(SaturatingCounter_82_reset),
    .io_enable(SaturatingCounter_82_io_enable),
    .io_value(SaturatingCounter_82_io_value)
  );
  SaturatingCounter SaturatingCounter_83 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_83_clock),
    .reset(SaturatingCounter_83_reset),
    .io_enable(SaturatingCounter_83_io_enable),
    .io_value(SaturatingCounter_83_io_value)
  );
  SaturatingCounter SaturatingCounter_84 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_84_clock),
    .reset(SaturatingCounter_84_reset),
    .io_enable(SaturatingCounter_84_io_enable),
    .io_value(SaturatingCounter_84_io_value)
  );
  SaturatingCounter SaturatingCounter_85 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_85_clock),
    .reset(SaturatingCounter_85_reset),
    .io_enable(SaturatingCounter_85_io_enable),
    .io_value(SaturatingCounter_85_io_value)
  );
  SaturatingCounter SaturatingCounter_86 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_86_clock),
    .reset(SaturatingCounter_86_reset),
    .io_enable(SaturatingCounter_86_io_enable),
    .io_value(SaturatingCounter_86_io_value)
  );
  SaturatingCounter SaturatingCounter_87 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_87_clock),
    .reset(SaturatingCounter_87_reset),
    .io_enable(SaturatingCounter_87_io_enable),
    .io_value(SaturatingCounter_87_io_value)
  );
  SaturatingCounter SaturatingCounter_88 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_88_clock),
    .reset(SaturatingCounter_88_reset),
    .io_enable(SaturatingCounter_88_io_enable),
    .io_value(SaturatingCounter_88_io_value)
  );
  SaturatingCounter SaturatingCounter_89 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_89_clock),
    .reset(SaturatingCounter_89_reset),
    .io_enable(SaturatingCounter_89_io_enable),
    .io_value(SaturatingCounter_89_io_value)
  );
  SaturatingCounter SaturatingCounter_90 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_90_clock),
    .reset(SaturatingCounter_90_reset),
    .io_enable(SaturatingCounter_90_io_enable),
    .io_value(SaturatingCounter_90_io_value)
  );
  SaturatingCounter SaturatingCounter_91 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_91_clock),
    .reset(SaturatingCounter_91_reset),
    .io_enable(SaturatingCounter_91_io_enable),
    .io_value(SaturatingCounter_91_io_value)
  );
  SaturatingCounter SaturatingCounter_92 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_92_clock),
    .reset(SaturatingCounter_92_reset),
    .io_enable(SaturatingCounter_92_io_enable),
    .io_value(SaturatingCounter_92_io_value)
  );
  SaturatingCounter SaturatingCounter_93 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_93_clock),
    .reset(SaturatingCounter_93_reset),
    .io_enable(SaturatingCounter_93_io_enable),
    .io_value(SaturatingCounter_93_io_value)
  );
  SaturatingCounter SaturatingCounter_94 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_94_clock),
    .reset(SaturatingCounter_94_reset),
    .io_enable(SaturatingCounter_94_io_enable),
    .io_value(SaturatingCounter_94_io_value)
  );
  SaturatingCounter SaturatingCounter_95 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_95_clock),
    .reset(SaturatingCounter_95_reset),
    .io_enable(SaturatingCounter_95_io_enable),
    .io_value(SaturatingCounter_95_io_value)
  );
  SaturatingCounter SaturatingCounter_96 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_96_clock),
    .reset(SaturatingCounter_96_reset),
    .io_enable(SaturatingCounter_96_io_enable),
    .io_value(SaturatingCounter_96_io_value)
  );
  SaturatingCounter SaturatingCounter_97 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_97_clock),
    .reset(SaturatingCounter_97_reset),
    .io_enable(SaturatingCounter_97_io_enable),
    .io_value(SaturatingCounter_97_io_value)
  );
  SaturatingCounter SaturatingCounter_98 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_98_clock),
    .reset(SaturatingCounter_98_reset),
    .io_enable(SaturatingCounter_98_io_enable),
    .io_value(SaturatingCounter_98_io_value)
  );
  SaturatingCounter SaturatingCounter_99 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_99_clock),
    .reset(SaturatingCounter_99_reset),
    .io_enable(SaturatingCounter_99_io_enable),
    .io_value(SaturatingCounter_99_io_value)
  );
  SaturatingCounter SaturatingCounter_100 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_100_clock),
    .reset(SaturatingCounter_100_reset),
    .io_enable(SaturatingCounter_100_io_enable),
    .io_value(SaturatingCounter_100_io_value)
  );
  SaturatingCounter SaturatingCounter_101 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_101_clock),
    .reset(SaturatingCounter_101_reset),
    .io_enable(SaturatingCounter_101_io_enable),
    .io_value(SaturatingCounter_101_io_value)
  );
  SaturatingCounter SaturatingCounter_102 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_102_clock),
    .reset(SaturatingCounter_102_reset),
    .io_enable(SaturatingCounter_102_io_enable),
    .io_value(SaturatingCounter_102_io_value)
  );
  SaturatingCounter SaturatingCounter_103 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_103_clock),
    .reset(SaturatingCounter_103_reset),
    .io_enable(SaturatingCounter_103_io_enable),
    .io_value(SaturatingCounter_103_io_value)
  );
  SaturatingCounter SaturatingCounter_104 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_104_clock),
    .reset(SaturatingCounter_104_reset),
    .io_enable(SaturatingCounter_104_io_enable),
    .io_value(SaturatingCounter_104_io_value)
  );
  SaturatingCounter SaturatingCounter_105 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_105_clock),
    .reset(SaturatingCounter_105_reset),
    .io_enable(SaturatingCounter_105_io_enable),
    .io_value(SaturatingCounter_105_io_value)
  );
  SaturatingCounter SaturatingCounter_106 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_106_clock),
    .reset(SaturatingCounter_106_reset),
    .io_enable(SaturatingCounter_106_io_enable),
    .io_value(SaturatingCounter_106_io_value)
  );
  SaturatingCounter SaturatingCounter_107 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_107_clock),
    .reset(SaturatingCounter_107_reset),
    .io_enable(SaturatingCounter_107_io_enable),
    .io_value(SaturatingCounter_107_io_value)
  );
  SaturatingCounter SaturatingCounter_108 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_108_clock),
    .reset(SaturatingCounter_108_reset),
    .io_enable(SaturatingCounter_108_io_enable),
    .io_value(SaturatingCounter_108_io_value)
  );
  SaturatingCounter SaturatingCounter_109 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_109_clock),
    .reset(SaturatingCounter_109_reset),
    .io_enable(SaturatingCounter_109_io_enable),
    .io_value(SaturatingCounter_109_io_value)
  );
  SaturatingCounter SaturatingCounter_110 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_110_clock),
    .reset(SaturatingCounter_110_reset),
    .io_enable(SaturatingCounter_110_io_enable),
    .io_value(SaturatingCounter_110_io_value)
  );
  SaturatingCounter SaturatingCounter_111 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_111_clock),
    .reset(SaturatingCounter_111_reset),
    .io_enable(SaturatingCounter_111_io_enable),
    .io_value(SaturatingCounter_111_io_value)
  );
  SaturatingCounter SaturatingCounter_112 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_112_clock),
    .reset(SaturatingCounter_112_reset),
    .io_enable(SaturatingCounter_112_io_enable),
    .io_value(SaturatingCounter_112_io_value)
  );
  SaturatingCounter SaturatingCounter_113 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_113_clock),
    .reset(SaturatingCounter_113_reset),
    .io_enable(SaturatingCounter_113_io_enable),
    .io_value(SaturatingCounter_113_io_value)
  );
  SaturatingCounter SaturatingCounter_114 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_114_clock),
    .reset(SaturatingCounter_114_reset),
    .io_enable(SaturatingCounter_114_io_enable),
    .io_value(SaturatingCounter_114_io_value)
  );
  SaturatingCounter SaturatingCounter_115 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_115_clock),
    .reset(SaturatingCounter_115_reset),
    .io_enable(SaturatingCounter_115_io_enable),
    .io_value(SaturatingCounter_115_io_value)
  );
  SaturatingCounter SaturatingCounter_116 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_116_clock),
    .reset(SaturatingCounter_116_reset),
    .io_enable(SaturatingCounter_116_io_enable),
    .io_value(SaturatingCounter_116_io_value)
  );
  SaturatingCounter SaturatingCounter_117 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_117_clock),
    .reset(SaturatingCounter_117_reset),
    .io_enable(SaturatingCounter_117_io_enable),
    .io_value(SaturatingCounter_117_io_value)
  );
  SaturatingCounter SaturatingCounter_118 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_118_clock),
    .reset(SaturatingCounter_118_reset),
    .io_enable(SaturatingCounter_118_io_enable),
    .io_value(SaturatingCounter_118_io_value)
  );
  SaturatingCounter SaturatingCounter_119 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_119_clock),
    .reset(SaturatingCounter_119_reset),
    .io_enable(SaturatingCounter_119_io_enable),
    .io_value(SaturatingCounter_119_io_value)
  );
  SaturatingCounter SaturatingCounter_120 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_120_clock),
    .reset(SaturatingCounter_120_reset),
    .io_enable(SaturatingCounter_120_io_enable),
    .io_value(SaturatingCounter_120_io_value)
  );
  SaturatingCounter SaturatingCounter_121 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_121_clock),
    .reset(SaturatingCounter_121_reset),
    .io_enable(SaturatingCounter_121_io_enable),
    .io_value(SaturatingCounter_121_io_value)
  );
  SaturatingCounter SaturatingCounter_122 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_122_clock),
    .reset(SaturatingCounter_122_reset),
    .io_enable(SaturatingCounter_122_io_enable),
    .io_value(SaturatingCounter_122_io_value)
  );
  SaturatingCounter SaturatingCounter_123 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_123_clock),
    .reset(SaturatingCounter_123_reset),
    .io_enable(SaturatingCounter_123_io_enable),
    .io_value(SaturatingCounter_123_io_value)
  );
  SaturatingCounter SaturatingCounter_124 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_124_clock),
    .reset(SaturatingCounter_124_reset),
    .io_enable(SaturatingCounter_124_io_enable),
    .io_value(SaturatingCounter_124_io_value)
  );
  SaturatingCounter SaturatingCounter_125 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_125_clock),
    .reset(SaturatingCounter_125_reset),
    .io_enable(SaturatingCounter_125_io_enable),
    .io_value(SaturatingCounter_125_io_value)
  );
  SaturatingCounter SaturatingCounter_126 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_126_clock),
    .reset(SaturatingCounter_126_reset),
    .io_enable(SaturatingCounter_126_io_enable),
    .io_value(SaturatingCounter_126_io_value)
  );
  SaturatingCounter SaturatingCounter_127 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_127_clock),
    .reset(SaturatingCounter_127_reset),
    .io_enable(SaturatingCounter_127_io_enable),
    .io_value(SaturatingCounter_127_io_value)
  );
  SaturatingCounter SaturatingCounter_128 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_128_clock),
    .reset(SaturatingCounter_128_reset),
    .io_enable(SaturatingCounter_128_io_enable),
    .io_value(SaturatingCounter_128_io_value)
  );
  SaturatingCounter SaturatingCounter_129 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_129_clock),
    .reset(SaturatingCounter_129_reset),
    .io_enable(SaturatingCounter_129_io_enable),
    .io_value(SaturatingCounter_129_io_value)
  );
  SaturatingCounter SaturatingCounter_130 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_130_clock),
    .reset(SaturatingCounter_130_reset),
    .io_enable(SaturatingCounter_130_io_enable),
    .io_value(SaturatingCounter_130_io_value)
  );
  SaturatingCounter SaturatingCounter_131 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_131_clock),
    .reset(SaturatingCounter_131_reset),
    .io_enable(SaturatingCounter_131_io_enable),
    .io_value(SaturatingCounter_131_io_value)
  );
  SaturatingCounter SaturatingCounter_132 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_132_clock),
    .reset(SaturatingCounter_132_reset),
    .io_enable(SaturatingCounter_132_io_enable),
    .io_value(SaturatingCounter_132_io_value)
  );
  SaturatingCounter SaturatingCounter_133 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_133_clock),
    .reset(SaturatingCounter_133_reset),
    .io_enable(SaturatingCounter_133_io_enable),
    .io_value(SaturatingCounter_133_io_value)
  );
  SaturatingCounter SaturatingCounter_134 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_134_clock),
    .reset(SaturatingCounter_134_reset),
    .io_enable(SaturatingCounter_134_io_enable),
    .io_value(SaturatingCounter_134_io_value)
  );
  SaturatingCounter SaturatingCounter_135 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_135_clock),
    .reset(SaturatingCounter_135_reset),
    .io_enable(SaturatingCounter_135_io_enable),
    .io_value(SaturatingCounter_135_io_value)
  );
  SaturatingCounter SaturatingCounter_136 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_136_clock),
    .reset(SaturatingCounter_136_reset),
    .io_enable(SaturatingCounter_136_io_enable),
    .io_value(SaturatingCounter_136_io_value)
  );
  SaturatingCounter SaturatingCounter_137 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_137_clock),
    .reset(SaturatingCounter_137_reset),
    .io_enable(SaturatingCounter_137_io_enable),
    .io_value(SaturatingCounter_137_io_value)
  );
  SaturatingCounter SaturatingCounter_138 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_138_clock),
    .reset(SaturatingCounter_138_reset),
    .io_enable(SaturatingCounter_138_io_enable),
    .io_value(SaturatingCounter_138_io_value)
  );
  SaturatingCounter SaturatingCounter_139 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_139_clock),
    .reset(SaturatingCounter_139_reset),
    .io_enable(SaturatingCounter_139_io_enable),
    .io_value(SaturatingCounter_139_io_value)
  );
  SaturatingCounter SaturatingCounter_140 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_140_clock),
    .reset(SaturatingCounter_140_reset),
    .io_enable(SaturatingCounter_140_io_enable),
    .io_value(SaturatingCounter_140_io_value)
  );
  SaturatingCounter SaturatingCounter_141 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_141_clock),
    .reset(SaturatingCounter_141_reset),
    .io_enable(SaturatingCounter_141_io_enable),
    .io_value(SaturatingCounter_141_io_value)
  );
  SaturatingCounter SaturatingCounter_142 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_142_clock),
    .reset(SaturatingCounter_142_reset),
    .io_enable(SaturatingCounter_142_io_enable),
    .io_value(SaturatingCounter_142_io_value)
  );
  SaturatingCounter SaturatingCounter_143 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_143_clock),
    .reset(SaturatingCounter_143_reset),
    .io_enable(SaturatingCounter_143_io_enable),
    .io_value(SaturatingCounter_143_io_value)
  );
  SaturatingCounter SaturatingCounter_144 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_144_clock),
    .reset(SaturatingCounter_144_reset),
    .io_enable(SaturatingCounter_144_io_enable),
    .io_value(SaturatingCounter_144_io_value)
  );
  SaturatingCounter SaturatingCounter_145 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_145_clock),
    .reset(SaturatingCounter_145_reset),
    .io_enable(SaturatingCounter_145_io_enable),
    .io_value(SaturatingCounter_145_io_value)
  );
  SaturatingCounter SaturatingCounter_146 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_146_clock),
    .reset(SaturatingCounter_146_reset),
    .io_enable(SaturatingCounter_146_io_enable),
    .io_value(SaturatingCounter_146_io_value)
  );
  SaturatingCounter SaturatingCounter_147 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_147_clock),
    .reset(SaturatingCounter_147_reset),
    .io_enable(SaturatingCounter_147_io_enable),
    .io_value(SaturatingCounter_147_io_value)
  );
  SaturatingCounter SaturatingCounter_148 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_148_clock),
    .reset(SaturatingCounter_148_reset),
    .io_enable(SaturatingCounter_148_io_enable),
    .io_value(SaturatingCounter_148_io_value)
  );
  SaturatingCounter SaturatingCounter_149 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_149_clock),
    .reset(SaturatingCounter_149_reset),
    .io_enable(SaturatingCounter_149_io_enable),
    .io_value(SaturatingCounter_149_io_value)
  );
  SaturatingCounter SaturatingCounter_150 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_150_clock),
    .reset(SaturatingCounter_150_reset),
    .io_enable(SaturatingCounter_150_io_enable),
    .io_value(SaturatingCounter_150_io_value)
  );
  SaturatingCounter SaturatingCounter_151 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_151_clock),
    .reset(SaturatingCounter_151_reset),
    .io_enable(SaturatingCounter_151_io_enable),
    .io_value(SaturatingCounter_151_io_value)
  );
  SaturatingCounter SaturatingCounter_152 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_152_clock),
    .reset(SaturatingCounter_152_reset),
    .io_enable(SaturatingCounter_152_io_enable),
    .io_value(SaturatingCounter_152_io_value)
  );
  SaturatingCounter SaturatingCounter_153 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_153_clock),
    .reset(SaturatingCounter_153_reset),
    .io_enable(SaturatingCounter_153_io_enable),
    .io_value(SaturatingCounter_153_io_value)
  );
  SaturatingCounter SaturatingCounter_154 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_154_clock),
    .reset(SaturatingCounter_154_reset),
    .io_enable(SaturatingCounter_154_io_enable),
    .io_value(SaturatingCounter_154_io_value)
  );
  SaturatingCounter SaturatingCounter_155 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_155_clock),
    .reset(SaturatingCounter_155_reset),
    .io_enable(SaturatingCounter_155_io_enable),
    .io_value(SaturatingCounter_155_io_value)
  );
  SaturatingCounter SaturatingCounter_156 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_156_clock),
    .reset(SaturatingCounter_156_reset),
    .io_enable(SaturatingCounter_156_io_enable),
    .io_value(SaturatingCounter_156_io_value)
  );
  SaturatingCounter SaturatingCounter_157 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_157_clock),
    .reset(SaturatingCounter_157_reset),
    .io_enable(SaturatingCounter_157_io_enable),
    .io_value(SaturatingCounter_157_io_value)
  );
  SaturatingCounter SaturatingCounter_158 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_158_clock),
    .reset(SaturatingCounter_158_reset),
    .io_enable(SaturatingCounter_158_io_enable),
    .io_value(SaturatingCounter_158_io_value)
  );
  SaturatingCounter SaturatingCounter_159 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_159_clock),
    .reset(SaturatingCounter_159_reset),
    .io_enable(SaturatingCounter_159_io_enable),
    .io_value(SaturatingCounter_159_io_value)
  );
  SaturatingCounter SaturatingCounter_160 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_160_clock),
    .reset(SaturatingCounter_160_reset),
    .io_enable(SaturatingCounter_160_io_enable),
    .io_value(SaturatingCounter_160_io_value)
  );
  SaturatingCounter SaturatingCounter_161 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_161_clock),
    .reset(SaturatingCounter_161_reset),
    .io_enable(SaturatingCounter_161_io_enable),
    .io_value(SaturatingCounter_161_io_value)
  );
  SaturatingCounter SaturatingCounter_162 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_162_clock),
    .reset(SaturatingCounter_162_reset),
    .io_enable(SaturatingCounter_162_io_enable),
    .io_value(SaturatingCounter_162_io_value)
  );
  SaturatingCounter SaturatingCounter_163 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_163_clock),
    .reset(SaturatingCounter_163_reset),
    .io_enable(SaturatingCounter_163_io_enable),
    .io_value(SaturatingCounter_163_io_value)
  );
  SaturatingCounter SaturatingCounter_164 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_164_clock),
    .reset(SaturatingCounter_164_reset),
    .io_enable(SaturatingCounter_164_io_enable),
    .io_value(SaturatingCounter_164_io_value)
  );
  SaturatingCounter SaturatingCounter_165 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_165_clock),
    .reset(SaturatingCounter_165_reset),
    .io_enable(SaturatingCounter_165_io_enable),
    .io_value(SaturatingCounter_165_io_value)
  );
  SaturatingCounter SaturatingCounter_166 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_166_clock),
    .reset(SaturatingCounter_166_reset),
    .io_enable(SaturatingCounter_166_io_enable),
    .io_value(SaturatingCounter_166_io_value)
  );
  SaturatingCounter SaturatingCounter_167 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_167_clock),
    .reset(SaturatingCounter_167_reset),
    .io_enable(SaturatingCounter_167_io_enable),
    .io_value(SaturatingCounter_167_io_value)
  );
  SaturatingCounter SaturatingCounter_168 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_168_clock),
    .reset(SaturatingCounter_168_reset),
    .io_enable(SaturatingCounter_168_io_enable),
    .io_value(SaturatingCounter_168_io_value)
  );
  SaturatingCounter SaturatingCounter_169 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_169_clock),
    .reset(SaturatingCounter_169_reset),
    .io_enable(SaturatingCounter_169_io_enable),
    .io_value(SaturatingCounter_169_io_value)
  );
  SaturatingCounter SaturatingCounter_170 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_170_clock),
    .reset(SaturatingCounter_170_reset),
    .io_enable(SaturatingCounter_170_io_enable),
    .io_value(SaturatingCounter_170_io_value)
  );
  SaturatingCounter SaturatingCounter_171 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_171_clock),
    .reset(SaturatingCounter_171_reset),
    .io_enable(SaturatingCounter_171_io_enable),
    .io_value(SaturatingCounter_171_io_value)
  );
  SaturatingCounter SaturatingCounter_172 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_172_clock),
    .reset(SaturatingCounter_172_reset),
    .io_enable(SaturatingCounter_172_io_enable),
    .io_value(SaturatingCounter_172_io_value)
  );
  SaturatingCounter SaturatingCounter_173 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_173_clock),
    .reset(SaturatingCounter_173_reset),
    .io_enable(SaturatingCounter_173_io_enable),
    .io_value(SaturatingCounter_173_io_value)
  );
  SaturatingCounter SaturatingCounter_174 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_174_clock),
    .reset(SaturatingCounter_174_reset),
    .io_enable(SaturatingCounter_174_io_enable),
    .io_value(SaturatingCounter_174_io_value)
  );
  SaturatingCounter SaturatingCounter_175 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_175_clock),
    .reset(SaturatingCounter_175_reset),
    .io_enable(SaturatingCounter_175_io_enable),
    .io_value(SaturatingCounter_175_io_value)
  );
  SaturatingCounter SaturatingCounter_176 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_176_clock),
    .reset(SaturatingCounter_176_reset),
    .io_enable(SaturatingCounter_176_io_enable),
    .io_value(SaturatingCounter_176_io_value)
  );
  SaturatingCounter SaturatingCounter_177 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_177_clock),
    .reset(SaturatingCounter_177_reset),
    .io_enable(SaturatingCounter_177_io_enable),
    .io_value(SaturatingCounter_177_io_value)
  );
  SaturatingCounter SaturatingCounter_178 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_178_clock),
    .reset(SaturatingCounter_178_reset),
    .io_enable(SaturatingCounter_178_io_enable),
    .io_value(SaturatingCounter_178_io_value)
  );
  SaturatingCounter SaturatingCounter_179 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_179_clock),
    .reset(SaturatingCounter_179_reset),
    .io_enable(SaturatingCounter_179_io_enable),
    .io_value(SaturatingCounter_179_io_value)
  );
  SaturatingCounter SaturatingCounter_180 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_180_clock),
    .reset(SaturatingCounter_180_reset),
    .io_enable(SaturatingCounter_180_io_enable),
    .io_value(SaturatingCounter_180_io_value)
  );
  SaturatingCounter SaturatingCounter_181 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_181_clock),
    .reset(SaturatingCounter_181_reset),
    .io_enable(SaturatingCounter_181_io_enable),
    .io_value(SaturatingCounter_181_io_value)
  );
  SaturatingCounter SaturatingCounter_182 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_182_clock),
    .reset(SaturatingCounter_182_reset),
    .io_enable(SaturatingCounter_182_io_enable),
    .io_value(SaturatingCounter_182_io_value)
  );
  SaturatingCounter SaturatingCounter_183 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_183_clock),
    .reset(SaturatingCounter_183_reset),
    .io_enable(SaturatingCounter_183_io_enable),
    .io_value(SaturatingCounter_183_io_value)
  );
  SaturatingCounter SaturatingCounter_184 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_184_clock),
    .reset(SaturatingCounter_184_reset),
    .io_enable(SaturatingCounter_184_io_enable),
    .io_value(SaturatingCounter_184_io_value)
  );
  SaturatingCounter SaturatingCounter_185 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_185_clock),
    .reset(SaturatingCounter_185_reset),
    .io_enable(SaturatingCounter_185_io_enable),
    .io_value(SaturatingCounter_185_io_value)
  );
  SaturatingCounter SaturatingCounter_186 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_186_clock),
    .reset(SaturatingCounter_186_reset),
    .io_enable(SaturatingCounter_186_io_enable),
    .io_value(SaturatingCounter_186_io_value)
  );
  SaturatingCounter SaturatingCounter_187 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_187_clock),
    .reset(SaturatingCounter_187_reset),
    .io_enable(SaturatingCounter_187_io_enable),
    .io_value(SaturatingCounter_187_io_value)
  );
  SaturatingCounter SaturatingCounter_188 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_188_clock),
    .reset(SaturatingCounter_188_reset),
    .io_enable(SaturatingCounter_188_io_enable),
    .io_value(SaturatingCounter_188_io_value)
  );
  SaturatingCounter SaturatingCounter_189 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_189_clock),
    .reset(SaturatingCounter_189_reset),
    .io_enable(SaturatingCounter_189_io_enable),
    .io_value(SaturatingCounter_189_io_value)
  );
  SaturatingCounter SaturatingCounter_190 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_190_clock),
    .reset(SaturatingCounter_190_reset),
    .io_enable(SaturatingCounter_190_io_enable),
    .io_value(SaturatingCounter_190_io_value)
  );
  SaturatingCounter SaturatingCounter_191 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_191_clock),
    .reset(SaturatingCounter_191_reset),
    .io_enable(SaturatingCounter_191_io_enable),
    .io_value(SaturatingCounter_191_io_value)
  );
  SaturatingCounter SaturatingCounter_192 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_192_clock),
    .reset(SaturatingCounter_192_reset),
    .io_enable(SaturatingCounter_192_io_enable),
    .io_value(SaturatingCounter_192_io_value)
  );
  SaturatingCounter SaturatingCounter_193 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_193_clock),
    .reset(SaturatingCounter_193_reset),
    .io_enable(SaturatingCounter_193_io_enable),
    .io_value(SaturatingCounter_193_io_value)
  );
  SaturatingCounter SaturatingCounter_194 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_194_clock),
    .reset(SaturatingCounter_194_reset),
    .io_enable(SaturatingCounter_194_io_enable),
    .io_value(SaturatingCounter_194_io_value)
  );
  SaturatingCounter SaturatingCounter_195 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_195_clock),
    .reset(SaturatingCounter_195_reset),
    .io_enable(SaturatingCounter_195_io_enable),
    .io_value(SaturatingCounter_195_io_value)
  );
  SaturatingCounter SaturatingCounter_196 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_196_clock),
    .reset(SaturatingCounter_196_reset),
    .io_enable(SaturatingCounter_196_io_enable),
    .io_value(SaturatingCounter_196_io_value)
  );
  SaturatingCounter SaturatingCounter_197 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_197_clock),
    .reset(SaturatingCounter_197_reset),
    .io_enable(SaturatingCounter_197_io_enable),
    .io_value(SaturatingCounter_197_io_value)
  );
  SaturatingCounter SaturatingCounter_198 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_198_clock),
    .reset(SaturatingCounter_198_reset),
    .io_enable(SaturatingCounter_198_io_enable),
    .io_value(SaturatingCounter_198_io_value)
  );
  SaturatingCounter SaturatingCounter_199 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_199_clock),
    .reset(SaturatingCounter_199_reset),
    .io_enable(SaturatingCounter_199_io_enable),
    .io_value(SaturatingCounter_199_io_value)
  );
  SaturatingCounter SaturatingCounter_200 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_200_clock),
    .reset(SaturatingCounter_200_reset),
    .io_enable(SaturatingCounter_200_io_enable),
    .io_value(SaturatingCounter_200_io_value)
  );
  SaturatingCounter SaturatingCounter_201 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_201_clock),
    .reset(SaturatingCounter_201_reset),
    .io_enable(SaturatingCounter_201_io_enable),
    .io_value(SaturatingCounter_201_io_value)
  );
  SaturatingCounter SaturatingCounter_202 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_202_clock),
    .reset(SaturatingCounter_202_reset),
    .io_enable(SaturatingCounter_202_io_enable),
    .io_value(SaturatingCounter_202_io_value)
  );
  SaturatingCounter SaturatingCounter_203 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_203_clock),
    .reset(SaturatingCounter_203_reset),
    .io_enable(SaturatingCounter_203_io_enable),
    .io_value(SaturatingCounter_203_io_value)
  );
  SaturatingCounter SaturatingCounter_204 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_204_clock),
    .reset(SaturatingCounter_204_reset),
    .io_enable(SaturatingCounter_204_io_enable),
    .io_value(SaturatingCounter_204_io_value)
  );
  SaturatingCounter SaturatingCounter_205 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_205_clock),
    .reset(SaturatingCounter_205_reset),
    .io_enable(SaturatingCounter_205_io_enable),
    .io_value(SaturatingCounter_205_io_value)
  );
  SaturatingCounter SaturatingCounter_206 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_206_clock),
    .reset(SaturatingCounter_206_reset),
    .io_enable(SaturatingCounter_206_io_enable),
    .io_value(SaturatingCounter_206_io_value)
  );
  SaturatingCounter SaturatingCounter_207 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_207_clock),
    .reset(SaturatingCounter_207_reset),
    .io_enable(SaturatingCounter_207_io_enable),
    .io_value(SaturatingCounter_207_io_value)
  );
  SaturatingCounter SaturatingCounter_208 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_208_clock),
    .reset(SaturatingCounter_208_reset),
    .io_enable(SaturatingCounter_208_io_enable),
    .io_value(SaturatingCounter_208_io_value)
  );
  SaturatingCounter SaturatingCounter_209 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_209_clock),
    .reset(SaturatingCounter_209_reset),
    .io_enable(SaturatingCounter_209_io_enable),
    .io_value(SaturatingCounter_209_io_value)
  );
  SaturatingCounter SaturatingCounter_210 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_210_clock),
    .reset(SaturatingCounter_210_reset),
    .io_enable(SaturatingCounter_210_io_enable),
    .io_value(SaturatingCounter_210_io_value)
  );
  SaturatingCounter SaturatingCounter_211 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_211_clock),
    .reset(SaturatingCounter_211_reset),
    .io_enable(SaturatingCounter_211_io_enable),
    .io_value(SaturatingCounter_211_io_value)
  );
  SaturatingCounter SaturatingCounter_212 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_212_clock),
    .reset(SaturatingCounter_212_reset),
    .io_enable(SaturatingCounter_212_io_enable),
    .io_value(SaturatingCounter_212_io_value)
  );
  SaturatingCounter SaturatingCounter_213 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_213_clock),
    .reset(SaturatingCounter_213_reset),
    .io_enable(SaturatingCounter_213_io_enable),
    .io_value(SaturatingCounter_213_io_value)
  );
  SaturatingCounter SaturatingCounter_214 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_214_clock),
    .reset(SaturatingCounter_214_reset),
    .io_enable(SaturatingCounter_214_io_enable),
    .io_value(SaturatingCounter_214_io_value)
  );
  SaturatingCounter SaturatingCounter_215 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_215_clock),
    .reset(SaturatingCounter_215_reset),
    .io_enable(SaturatingCounter_215_io_enable),
    .io_value(SaturatingCounter_215_io_value)
  );
  SaturatingCounter SaturatingCounter_216 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_216_clock),
    .reset(SaturatingCounter_216_reset),
    .io_enable(SaturatingCounter_216_io_enable),
    .io_value(SaturatingCounter_216_io_value)
  );
  SaturatingCounter SaturatingCounter_217 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_217_clock),
    .reset(SaturatingCounter_217_reset),
    .io_enable(SaturatingCounter_217_io_enable),
    .io_value(SaturatingCounter_217_io_value)
  );
  SaturatingCounter SaturatingCounter_218 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_218_clock),
    .reset(SaturatingCounter_218_reset),
    .io_enable(SaturatingCounter_218_io_enable),
    .io_value(SaturatingCounter_218_io_value)
  );
  SaturatingCounter SaturatingCounter_219 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_219_clock),
    .reset(SaturatingCounter_219_reset),
    .io_enable(SaturatingCounter_219_io_enable),
    .io_value(SaturatingCounter_219_io_value)
  );
  SaturatingCounter SaturatingCounter_220 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_220_clock),
    .reset(SaturatingCounter_220_reset),
    .io_enable(SaturatingCounter_220_io_enable),
    .io_value(SaturatingCounter_220_io_value)
  );
  SaturatingCounter SaturatingCounter_221 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_221_clock),
    .reset(SaturatingCounter_221_reset),
    .io_enable(SaturatingCounter_221_io_enable),
    .io_value(SaturatingCounter_221_io_value)
  );
  SaturatingCounter SaturatingCounter_222 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_222_clock),
    .reset(SaturatingCounter_222_reset),
    .io_enable(SaturatingCounter_222_io_enable),
    .io_value(SaturatingCounter_222_io_value)
  );
  SaturatingCounter SaturatingCounter_223 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_223_clock),
    .reset(SaturatingCounter_223_reset),
    .io_enable(SaturatingCounter_223_io_enable),
    .io_value(SaturatingCounter_223_io_value)
  );
  SaturatingCounter SaturatingCounter_224 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_224_clock),
    .reset(SaturatingCounter_224_reset),
    .io_enable(SaturatingCounter_224_io_enable),
    .io_value(SaturatingCounter_224_io_value)
  );
  SaturatingCounter SaturatingCounter_225 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_225_clock),
    .reset(SaturatingCounter_225_reset),
    .io_enable(SaturatingCounter_225_io_enable),
    .io_value(SaturatingCounter_225_io_value)
  );
  SaturatingCounter SaturatingCounter_226 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_226_clock),
    .reset(SaturatingCounter_226_reset),
    .io_enable(SaturatingCounter_226_io_enable),
    .io_value(SaturatingCounter_226_io_value)
  );
  SaturatingCounter SaturatingCounter_227 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_227_clock),
    .reset(SaturatingCounter_227_reset),
    .io_enable(SaturatingCounter_227_io_enable),
    .io_value(SaturatingCounter_227_io_value)
  );
  SaturatingCounter SaturatingCounter_228 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_228_clock),
    .reset(SaturatingCounter_228_reset),
    .io_enable(SaturatingCounter_228_io_enable),
    .io_value(SaturatingCounter_228_io_value)
  );
  SaturatingCounter SaturatingCounter_229 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_229_clock),
    .reset(SaturatingCounter_229_reset),
    .io_enable(SaturatingCounter_229_io_enable),
    .io_value(SaturatingCounter_229_io_value)
  );
  SaturatingCounter SaturatingCounter_230 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_230_clock),
    .reset(SaturatingCounter_230_reset),
    .io_enable(SaturatingCounter_230_io_enable),
    .io_value(SaturatingCounter_230_io_value)
  );
  SaturatingCounter SaturatingCounter_231 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_231_clock),
    .reset(SaturatingCounter_231_reset),
    .io_enable(SaturatingCounter_231_io_enable),
    .io_value(SaturatingCounter_231_io_value)
  );
  SaturatingCounter SaturatingCounter_232 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_232_clock),
    .reset(SaturatingCounter_232_reset),
    .io_enable(SaturatingCounter_232_io_enable),
    .io_value(SaturatingCounter_232_io_value)
  );
  SaturatingCounter SaturatingCounter_233 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_233_clock),
    .reset(SaturatingCounter_233_reset),
    .io_enable(SaturatingCounter_233_io_enable),
    .io_value(SaturatingCounter_233_io_value)
  );
  SaturatingCounter SaturatingCounter_234 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_234_clock),
    .reset(SaturatingCounter_234_reset),
    .io_enable(SaturatingCounter_234_io_enable),
    .io_value(SaturatingCounter_234_io_value)
  );
  SaturatingCounter SaturatingCounter_235 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_235_clock),
    .reset(SaturatingCounter_235_reset),
    .io_enable(SaturatingCounter_235_io_enable),
    .io_value(SaturatingCounter_235_io_value)
  );
  SaturatingCounter SaturatingCounter_236 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_236_clock),
    .reset(SaturatingCounter_236_reset),
    .io_enable(SaturatingCounter_236_io_enable),
    .io_value(SaturatingCounter_236_io_value)
  );
  SaturatingCounter SaturatingCounter_237 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_237_clock),
    .reset(SaturatingCounter_237_reset),
    .io_enable(SaturatingCounter_237_io_enable),
    .io_value(SaturatingCounter_237_io_value)
  );
  SaturatingCounter SaturatingCounter_238 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_238_clock),
    .reset(SaturatingCounter_238_reset),
    .io_enable(SaturatingCounter_238_io_enable),
    .io_value(SaturatingCounter_238_io_value)
  );
  SaturatingCounter SaturatingCounter_239 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_239_clock),
    .reset(SaturatingCounter_239_reset),
    .io_enable(SaturatingCounter_239_io_enable),
    .io_value(SaturatingCounter_239_io_value)
  );
  SaturatingCounter SaturatingCounter_240 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_240_clock),
    .reset(SaturatingCounter_240_reset),
    .io_enable(SaturatingCounter_240_io_enable),
    .io_value(SaturatingCounter_240_io_value)
  );
  SaturatingCounter SaturatingCounter_241 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_241_clock),
    .reset(SaturatingCounter_241_reset),
    .io_enable(SaturatingCounter_241_io_enable),
    .io_value(SaturatingCounter_241_io_value)
  );
  SaturatingCounter SaturatingCounter_242 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_242_clock),
    .reset(SaturatingCounter_242_reset),
    .io_enable(SaturatingCounter_242_io_enable),
    .io_value(SaturatingCounter_242_io_value)
  );
  SaturatingCounter SaturatingCounter_243 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_243_clock),
    .reset(SaturatingCounter_243_reset),
    .io_enable(SaturatingCounter_243_io_enable),
    .io_value(SaturatingCounter_243_io_value)
  );
  SaturatingCounter SaturatingCounter_244 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_244_clock),
    .reset(SaturatingCounter_244_reset),
    .io_enable(SaturatingCounter_244_io_enable),
    .io_value(SaturatingCounter_244_io_value)
  );
  SaturatingCounter SaturatingCounter_245 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_245_clock),
    .reset(SaturatingCounter_245_reset),
    .io_enable(SaturatingCounter_245_io_enable),
    .io_value(SaturatingCounter_245_io_value)
  );
  SaturatingCounter SaturatingCounter_246 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_246_clock),
    .reset(SaturatingCounter_246_reset),
    .io_enable(SaturatingCounter_246_io_enable),
    .io_value(SaturatingCounter_246_io_value)
  );
  SaturatingCounter SaturatingCounter_247 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_247_clock),
    .reset(SaturatingCounter_247_reset),
    .io_enable(SaturatingCounter_247_io_enable),
    .io_value(SaturatingCounter_247_io_value)
  );
  SaturatingCounter SaturatingCounter_248 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_248_clock),
    .reset(SaturatingCounter_248_reset),
    .io_enable(SaturatingCounter_248_io_enable),
    .io_value(SaturatingCounter_248_io_value)
  );
  SaturatingCounter SaturatingCounter_249 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_249_clock),
    .reset(SaturatingCounter_249_reset),
    .io_enable(SaturatingCounter_249_io_enable),
    .io_value(SaturatingCounter_249_io_value)
  );
  SaturatingCounter SaturatingCounter_250 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_250_clock),
    .reset(SaturatingCounter_250_reset),
    .io_enable(SaturatingCounter_250_io_enable),
    .io_value(SaturatingCounter_250_io_value)
  );
  SaturatingCounter SaturatingCounter_251 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_251_clock),
    .reset(SaturatingCounter_251_reset),
    .io_enable(SaturatingCounter_251_io_enable),
    .io_value(SaturatingCounter_251_io_value)
  );
  SaturatingCounter SaturatingCounter_252 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_252_clock),
    .reset(SaturatingCounter_252_reset),
    .io_enable(SaturatingCounter_252_io_enable),
    .io_value(SaturatingCounter_252_io_value)
  );
  SaturatingCounter SaturatingCounter_253 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_253_clock),
    .reset(SaturatingCounter_253_reset),
    .io_enable(SaturatingCounter_253_io_enable),
    .io_value(SaturatingCounter_253_io_value)
  );
  SaturatingCounter SaturatingCounter_254 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_254_clock),
    .reset(SaturatingCounter_254_reset),
    .io_enable(SaturatingCounter_254_io_enable),
    .io_value(SaturatingCounter_254_io_value)
  );
  SaturatingCounter SaturatingCounter_255 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_255_clock),
    .reset(SaturatingCounter_255_reset),
    .io_enable(SaturatingCounter_255_io_enable),
    .io_value(SaturatingCounter_255_io_value)
  );
  SaturatingCounter SaturatingCounter_256 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_256_clock),
    .reset(SaturatingCounter_256_reset),
    .io_enable(SaturatingCounter_256_io_enable),
    .io_value(SaturatingCounter_256_io_value)
  );
  SaturatingCounter SaturatingCounter_257 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_257_clock),
    .reset(SaturatingCounter_257_reset),
    .io_enable(SaturatingCounter_257_io_enable),
    .io_value(SaturatingCounter_257_io_value)
  );
  SaturatingCounter SaturatingCounter_258 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_258_clock),
    .reset(SaturatingCounter_258_reset),
    .io_enable(SaturatingCounter_258_io_enable),
    .io_value(SaturatingCounter_258_io_value)
  );
  SaturatingCounter SaturatingCounter_259 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_259_clock),
    .reset(SaturatingCounter_259_reset),
    .io_enable(SaturatingCounter_259_io_enable),
    .io_value(SaturatingCounter_259_io_value)
  );
  SaturatingCounter SaturatingCounter_260 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_260_clock),
    .reset(SaturatingCounter_260_reset),
    .io_enable(SaturatingCounter_260_io_enable),
    .io_value(SaturatingCounter_260_io_value)
  );
  SaturatingCounter SaturatingCounter_261 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_261_clock),
    .reset(SaturatingCounter_261_reset),
    .io_enable(SaturatingCounter_261_io_enable),
    .io_value(SaturatingCounter_261_io_value)
  );
  SaturatingCounter SaturatingCounter_262 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_262_clock),
    .reset(SaturatingCounter_262_reset),
    .io_enable(SaturatingCounter_262_io_enable),
    .io_value(SaturatingCounter_262_io_value)
  );
  SaturatingCounter SaturatingCounter_263 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_263_clock),
    .reset(SaturatingCounter_263_reset),
    .io_enable(SaturatingCounter_263_io_enable),
    .io_value(SaturatingCounter_263_io_value)
  );
  SaturatingCounter SaturatingCounter_264 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_264_clock),
    .reset(SaturatingCounter_264_reset),
    .io_enable(SaturatingCounter_264_io_enable),
    .io_value(SaturatingCounter_264_io_value)
  );
  SaturatingCounter SaturatingCounter_265 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_265_clock),
    .reset(SaturatingCounter_265_reset),
    .io_enable(SaturatingCounter_265_io_enable),
    .io_value(SaturatingCounter_265_io_value)
  );
  SaturatingCounter SaturatingCounter_266 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_266_clock),
    .reset(SaturatingCounter_266_reset),
    .io_enable(SaturatingCounter_266_io_enable),
    .io_value(SaturatingCounter_266_io_value)
  );
  SaturatingCounter SaturatingCounter_267 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_267_clock),
    .reset(SaturatingCounter_267_reset),
    .io_enable(SaturatingCounter_267_io_enable),
    .io_value(SaturatingCounter_267_io_value)
  );
  SaturatingCounter SaturatingCounter_268 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_268_clock),
    .reset(SaturatingCounter_268_reset),
    .io_enable(SaturatingCounter_268_io_enable),
    .io_value(SaturatingCounter_268_io_value)
  );
  SaturatingCounter SaturatingCounter_269 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_269_clock),
    .reset(SaturatingCounter_269_reset),
    .io_enable(SaturatingCounter_269_io_enable),
    .io_value(SaturatingCounter_269_io_value)
  );
  SaturatingCounter SaturatingCounter_270 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_270_clock),
    .reset(SaturatingCounter_270_reset),
    .io_enable(SaturatingCounter_270_io_enable),
    .io_value(SaturatingCounter_270_io_value)
  );
  SaturatingCounter SaturatingCounter_271 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_271_clock),
    .reset(SaturatingCounter_271_reset),
    .io_enable(SaturatingCounter_271_io_enable),
    .io_value(SaturatingCounter_271_io_value)
  );
  SaturatingCounter SaturatingCounter_272 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_272_clock),
    .reset(SaturatingCounter_272_reset),
    .io_enable(SaturatingCounter_272_io_enable),
    .io_value(SaturatingCounter_272_io_value)
  );
  SaturatingCounter SaturatingCounter_273 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_273_clock),
    .reset(SaturatingCounter_273_reset),
    .io_enable(SaturatingCounter_273_io_enable),
    .io_value(SaturatingCounter_273_io_value)
  );
  SaturatingCounter SaturatingCounter_274 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_274_clock),
    .reset(SaturatingCounter_274_reset),
    .io_enable(SaturatingCounter_274_io_enable),
    .io_value(SaturatingCounter_274_io_value)
  );
  SaturatingCounter SaturatingCounter_275 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_275_clock),
    .reset(SaturatingCounter_275_reset),
    .io_enable(SaturatingCounter_275_io_enable),
    .io_value(SaturatingCounter_275_io_value)
  );
  SaturatingCounter SaturatingCounter_276 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_276_clock),
    .reset(SaturatingCounter_276_reset),
    .io_enable(SaturatingCounter_276_io_enable),
    .io_value(SaturatingCounter_276_io_value)
  );
  SaturatingCounter SaturatingCounter_277 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_277_clock),
    .reset(SaturatingCounter_277_reset),
    .io_enable(SaturatingCounter_277_io_enable),
    .io_value(SaturatingCounter_277_io_value)
  );
  SaturatingCounter SaturatingCounter_278 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_278_clock),
    .reset(SaturatingCounter_278_reset),
    .io_enable(SaturatingCounter_278_io_enable),
    .io_value(SaturatingCounter_278_io_value)
  );
  SaturatingCounter SaturatingCounter_279 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_279_clock),
    .reset(SaturatingCounter_279_reset),
    .io_enable(SaturatingCounter_279_io_enable),
    .io_value(SaturatingCounter_279_io_value)
  );
  SaturatingCounter SaturatingCounter_280 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_280_clock),
    .reset(SaturatingCounter_280_reset),
    .io_enable(SaturatingCounter_280_io_enable),
    .io_value(SaturatingCounter_280_io_value)
  );
  SaturatingCounter SaturatingCounter_281 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_281_clock),
    .reset(SaturatingCounter_281_reset),
    .io_enable(SaturatingCounter_281_io_enable),
    .io_value(SaturatingCounter_281_io_value)
  );
  SaturatingCounter SaturatingCounter_282 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_282_clock),
    .reset(SaturatingCounter_282_reset),
    .io_enable(SaturatingCounter_282_io_enable),
    .io_value(SaturatingCounter_282_io_value)
  );
  SaturatingCounter SaturatingCounter_283 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_283_clock),
    .reset(SaturatingCounter_283_reset),
    .io_enable(SaturatingCounter_283_io_enable),
    .io_value(SaturatingCounter_283_io_value)
  );
  SaturatingCounter SaturatingCounter_284 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_284_clock),
    .reset(SaturatingCounter_284_reset),
    .io_enable(SaturatingCounter_284_io_enable),
    .io_value(SaturatingCounter_284_io_value)
  );
  SaturatingCounter SaturatingCounter_285 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_285_clock),
    .reset(SaturatingCounter_285_reset),
    .io_enable(SaturatingCounter_285_io_enable),
    .io_value(SaturatingCounter_285_io_value)
  );
  SaturatingCounter SaturatingCounter_286 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_286_clock),
    .reset(SaturatingCounter_286_reset),
    .io_enable(SaturatingCounter_286_io_enable),
    .io_value(SaturatingCounter_286_io_value)
  );
  SaturatingCounter SaturatingCounter_287 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_287_clock),
    .reset(SaturatingCounter_287_reset),
    .io_enable(SaturatingCounter_287_io_enable),
    .io_value(SaturatingCounter_287_io_value)
  );
  SaturatingCounter SaturatingCounter_288 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_288_clock),
    .reset(SaturatingCounter_288_reset),
    .io_enable(SaturatingCounter_288_io_enable),
    .io_value(SaturatingCounter_288_io_value)
  );
  SaturatingCounter SaturatingCounter_289 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_289_clock),
    .reset(SaturatingCounter_289_reset),
    .io_enable(SaturatingCounter_289_io_enable),
    .io_value(SaturatingCounter_289_io_value)
  );
  SaturatingCounter SaturatingCounter_290 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_290_clock),
    .reset(SaturatingCounter_290_reset),
    .io_enable(SaturatingCounter_290_io_enable),
    .io_value(SaturatingCounter_290_io_value)
  );
  SaturatingCounter SaturatingCounter_291 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_291_clock),
    .reset(SaturatingCounter_291_reset),
    .io_enable(SaturatingCounter_291_io_enable),
    .io_value(SaturatingCounter_291_io_value)
  );
  SaturatingCounter SaturatingCounter_292 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_292_clock),
    .reset(SaturatingCounter_292_reset),
    .io_enable(SaturatingCounter_292_io_enable),
    .io_value(SaturatingCounter_292_io_value)
  );
  SaturatingCounter SaturatingCounter_293 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_293_clock),
    .reset(SaturatingCounter_293_reset),
    .io_enable(SaturatingCounter_293_io_enable),
    .io_value(SaturatingCounter_293_io_value)
  );
  SaturatingCounter SaturatingCounter_294 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_294_clock),
    .reset(SaturatingCounter_294_reset),
    .io_enable(SaturatingCounter_294_io_enable),
    .io_value(SaturatingCounter_294_io_value)
  );
  SaturatingCounter SaturatingCounter_295 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_295_clock),
    .reset(SaturatingCounter_295_reset),
    .io_enable(SaturatingCounter_295_io_enable),
    .io_value(SaturatingCounter_295_io_value)
  );
  SaturatingCounter SaturatingCounter_296 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_296_clock),
    .reset(SaturatingCounter_296_reset),
    .io_enable(SaturatingCounter_296_io_enable),
    .io_value(SaturatingCounter_296_io_value)
  );
  SaturatingCounter SaturatingCounter_297 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_297_clock),
    .reset(SaturatingCounter_297_reset),
    .io_enable(SaturatingCounter_297_io_enable),
    .io_value(SaturatingCounter_297_io_value)
  );
  SaturatingCounter SaturatingCounter_298 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_298_clock),
    .reset(SaturatingCounter_298_reset),
    .io_enable(SaturatingCounter_298_io_enable),
    .io_value(SaturatingCounter_298_io_value)
  );
  SaturatingCounter SaturatingCounter_299 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_299_clock),
    .reset(SaturatingCounter_299_reset),
    .io_enable(SaturatingCounter_299_io_enable),
    .io_value(SaturatingCounter_299_io_value)
  );
  SaturatingCounter SaturatingCounter_300 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_300_clock),
    .reset(SaturatingCounter_300_reset),
    .io_enable(SaturatingCounter_300_io_enable),
    .io_value(SaturatingCounter_300_io_value)
  );
  SaturatingCounter SaturatingCounter_301 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_301_clock),
    .reset(SaturatingCounter_301_reset),
    .io_enable(SaturatingCounter_301_io_enable),
    .io_value(SaturatingCounter_301_io_value)
  );
  SaturatingCounter SaturatingCounter_302 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_302_clock),
    .reset(SaturatingCounter_302_reset),
    .io_enable(SaturatingCounter_302_io_enable),
    .io_value(SaturatingCounter_302_io_value)
  );
  SaturatingCounter SaturatingCounter_303 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_303_clock),
    .reset(SaturatingCounter_303_reset),
    .io_enable(SaturatingCounter_303_io_enable),
    .io_value(SaturatingCounter_303_io_value)
  );
  SaturatingCounter SaturatingCounter_304 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_304_clock),
    .reset(SaturatingCounter_304_reset),
    .io_enable(SaturatingCounter_304_io_enable),
    .io_value(SaturatingCounter_304_io_value)
  );
  SaturatingCounter SaturatingCounter_305 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_305_clock),
    .reset(SaturatingCounter_305_reset),
    .io_enable(SaturatingCounter_305_io_enable),
    .io_value(SaturatingCounter_305_io_value)
  );
  SaturatingCounter SaturatingCounter_306 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_306_clock),
    .reset(SaturatingCounter_306_reset),
    .io_enable(SaturatingCounter_306_io_enable),
    .io_value(SaturatingCounter_306_io_value)
  );
  SaturatingCounter SaturatingCounter_307 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_307_clock),
    .reset(SaturatingCounter_307_reset),
    .io_enable(SaturatingCounter_307_io_enable),
    .io_value(SaturatingCounter_307_io_value)
  );
  SaturatingCounter SaturatingCounter_308 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_308_clock),
    .reset(SaturatingCounter_308_reset),
    .io_enable(SaturatingCounter_308_io_enable),
    .io_value(SaturatingCounter_308_io_value)
  );
  SaturatingCounter SaturatingCounter_309 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_309_clock),
    .reset(SaturatingCounter_309_reset),
    .io_enable(SaturatingCounter_309_io_enable),
    .io_value(SaturatingCounter_309_io_value)
  );
  SaturatingCounter SaturatingCounter_310 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_310_clock),
    .reset(SaturatingCounter_310_reset),
    .io_enable(SaturatingCounter_310_io_enable),
    .io_value(SaturatingCounter_310_io_value)
  );
  SaturatingCounter SaturatingCounter_311 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_311_clock),
    .reset(SaturatingCounter_311_reset),
    .io_enable(SaturatingCounter_311_io_enable),
    .io_value(SaturatingCounter_311_io_value)
  );
  SaturatingCounter SaturatingCounter_312 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_312_clock),
    .reset(SaturatingCounter_312_reset),
    .io_enable(SaturatingCounter_312_io_enable),
    .io_value(SaturatingCounter_312_io_value)
  );
  SaturatingCounter SaturatingCounter_313 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_313_clock),
    .reset(SaturatingCounter_313_reset),
    .io_enable(SaturatingCounter_313_io_enable),
    .io_value(SaturatingCounter_313_io_value)
  );
  SaturatingCounter SaturatingCounter_314 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_314_clock),
    .reset(SaturatingCounter_314_reset),
    .io_enable(SaturatingCounter_314_io_enable),
    .io_value(SaturatingCounter_314_io_value)
  );
  SaturatingCounter SaturatingCounter_315 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_315_clock),
    .reset(SaturatingCounter_315_reset),
    .io_enable(SaturatingCounter_315_io_enable),
    .io_value(SaturatingCounter_315_io_value)
  );
  SaturatingCounter SaturatingCounter_316 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_316_clock),
    .reset(SaturatingCounter_316_reset),
    .io_enable(SaturatingCounter_316_io_enable),
    .io_value(SaturatingCounter_316_io_value)
  );
  SaturatingCounter SaturatingCounter_317 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_317_clock),
    .reset(SaturatingCounter_317_reset),
    .io_enable(SaturatingCounter_317_io_enable),
    .io_value(SaturatingCounter_317_io_value)
  );
  SaturatingCounter SaturatingCounter_318 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_318_clock),
    .reset(SaturatingCounter_318_reset),
    .io_enable(SaturatingCounter_318_io_enable),
    .io_value(SaturatingCounter_318_io_value)
  );
  SaturatingCounter SaturatingCounter_319 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_319_clock),
    .reset(SaturatingCounter_319_reset),
    .io_enable(SaturatingCounter_319_io_enable),
    .io_value(SaturatingCounter_319_io_value)
  );
  SaturatingCounter SaturatingCounter_320 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_320_clock),
    .reset(SaturatingCounter_320_reset),
    .io_enable(SaturatingCounter_320_io_enable),
    .io_value(SaturatingCounter_320_io_value)
  );
  SaturatingCounter SaturatingCounter_321 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_321_clock),
    .reset(SaturatingCounter_321_reset),
    .io_enable(SaturatingCounter_321_io_enable),
    .io_value(SaturatingCounter_321_io_value)
  );
  SaturatingCounter SaturatingCounter_322 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_322_clock),
    .reset(SaturatingCounter_322_reset),
    .io_enable(SaturatingCounter_322_io_enable),
    .io_value(SaturatingCounter_322_io_value)
  );
  SaturatingCounter SaturatingCounter_323 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_323_clock),
    .reset(SaturatingCounter_323_reset),
    .io_enable(SaturatingCounter_323_io_enable),
    .io_value(SaturatingCounter_323_io_value)
  );
  SaturatingCounter SaturatingCounter_324 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_324_clock),
    .reset(SaturatingCounter_324_reset),
    .io_enable(SaturatingCounter_324_io_enable),
    .io_value(SaturatingCounter_324_io_value)
  );
  SaturatingCounter SaturatingCounter_325 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_325_clock),
    .reset(SaturatingCounter_325_reset),
    .io_enable(SaturatingCounter_325_io_enable),
    .io_value(SaturatingCounter_325_io_value)
  );
  SaturatingCounter SaturatingCounter_326 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_326_clock),
    .reset(SaturatingCounter_326_reset),
    .io_enable(SaturatingCounter_326_io_enable),
    .io_value(SaturatingCounter_326_io_value)
  );
  SaturatingCounter SaturatingCounter_327 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_327_clock),
    .reset(SaturatingCounter_327_reset),
    .io_enable(SaturatingCounter_327_io_enable),
    .io_value(SaturatingCounter_327_io_value)
  );
  SaturatingCounter SaturatingCounter_328 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_328_clock),
    .reset(SaturatingCounter_328_reset),
    .io_enable(SaturatingCounter_328_io_enable),
    .io_value(SaturatingCounter_328_io_value)
  );
  SaturatingCounter SaturatingCounter_329 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_329_clock),
    .reset(SaturatingCounter_329_reset),
    .io_enable(SaturatingCounter_329_io_enable),
    .io_value(SaturatingCounter_329_io_value)
  );
  SaturatingCounter SaturatingCounter_330 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_330_clock),
    .reset(SaturatingCounter_330_reset),
    .io_enable(SaturatingCounter_330_io_enable),
    .io_value(SaturatingCounter_330_io_value)
  );
  SaturatingCounter SaturatingCounter_331 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_331_clock),
    .reset(SaturatingCounter_331_reset),
    .io_enable(SaturatingCounter_331_io_enable),
    .io_value(SaturatingCounter_331_io_value)
  );
  SaturatingCounter SaturatingCounter_332 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_332_clock),
    .reset(SaturatingCounter_332_reset),
    .io_enable(SaturatingCounter_332_io_enable),
    .io_value(SaturatingCounter_332_io_value)
  );
  SaturatingCounter SaturatingCounter_333 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_333_clock),
    .reset(SaturatingCounter_333_reset),
    .io_enable(SaturatingCounter_333_io_enable),
    .io_value(SaturatingCounter_333_io_value)
  );
  SaturatingCounter SaturatingCounter_334 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_334_clock),
    .reset(SaturatingCounter_334_reset),
    .io_enable(SaturatingCounter_334_io_enable),
    .io_value(SaturatingCounter_334_io_value)
  );
  SaturatingCounter SaturatingCounter_335 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_335_clock),
    .reset(SaturatingCounter_335_reset),
    .io_enable(SaturatingCounter_335_io_enable),
    .io_value(SaturatingCounter_335_io_value)
  );
  SaturatingCounter SaturatingCounter_336 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_336_clock),
    .reset(SaturatingCounter_336_reset),
    .io_enable(SaturatingCounter_336_io_enable),
    .io_value(SaturatingCounter_336_io_value)
  );
  SaturatingCounter SaturatingCounter_337 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_337_clock),
    .reset(SaturatingCounter_337_reset),
    .io_enable(SaturatingCounter_337_io_enable),
    .io_value(SaturatingCounter_337_io_value)
  );
  SaturatingCounter SaturatingCounter_338 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_338_clock),
    .reset(SaturatingCounter_338_reset),
    .io_enable(SaturatingCounter_338_io_enable),
    .io_value(SaturatingCounter_338_io_value)
  );
  SaturatingCounter SaturatingCounter_339 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_339_clock),
    .reset(SaturatingCounter_339_reset),
    .io_enable(SaturatingCounter_339_io_enable),
    .io_value(SaturatingCounter_339_io_value)
  );
  SaturatingCounter SaturatingCounter_340 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_340_clock),
    .reset(SaturatingCounter_340_reset),
    .io_enable(SaturatingCounter_340_io_enable),
    .io_value(SaturatingCounter_340_io_value)
  );
  SaturatingCounter SaturatingCounter_341 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_341_clock),
    .reset(SaturatingCounter_341_reset),
    .io_enable(SaturatingCounter_341_io_enable),
    .io_value(SaturatingCounter_341_io_value)
  );
  SaturatingCounter SaturatingCounter_342 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_342_clock),
    .reset(SaturatingCounter_342_reset),
    .io_enable(SaturatingCounter_342_io_enable),
    .io_value(SaturatingCounter_342_io_value)
  );
  SaturatingCounter SaturatingCounter_343 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_343_clock),
    .reset(SaturatingCounter_343_reset),
    .io_enable(SaturatingCounter_343_io_enable),
    .io_value(SaturatingCounter_343_io_value)
  );
  SaturatingCounter SaturatingCounter_344 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_344_clock),
    .reset(SaturatingCounter_344_reset),
    .io_enable(SaturatingCounter_344_io_enable),
    .io_value(SaturatingCounter_344_io_value)
  );
  SaturatingCounter SaturatingCounter_345 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_345_clock),
    .reset(SaturatingCounter_345_reset),
    .io_enable(SaturatingCounter_345_io_enable),
    .io_value(SaturatingCounter_345_io_value)
  );
  SaturatingCounter SaturatingCounter_346 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_346_clock),
    .reset(SaturatingCounter_346_reset),
    .io_enable(SaturatingCounter_346_io_enable),
    .io_value(SaturatingCounter_346_io_value)
  );
  SaturatingCounter SaturatingCounter_347 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_347_clock),
    .reset(SaturatingCounter_347_reset),
    .io_enable(SaturatingCounter_347_io_enable),
    .io_value(SaturatingCounter_347_io_value)
  );
  SaturatingCounter SaturatingCounter_348 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_348_clock),
    .reset(SaturatingCounter_348_reset),
    .io_enable(SaturatingCounter_348_io_enable),
    .io_value(SaturatingCounter_348_io_value)
  );
  SaturatingCounter SaturatingCounter_349 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_349_clock),
    .reset(SaturatingCounter_349_reset),
    .io_enable(SaturatingCounter_349_io_enable),
    .io_value(SaturatingCounter_349_io_value)
  );
  SaturatingCounter SaturatingCounter_350 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_350_clock),
    .reset(SaturatingCounter_350_reset),
    .io_enable(SaturatingCounter_350_io_enable),
    .io_value(SaturatingCounter_350_io_value)
  );
  SaturatingCounter SaturatingCounter_351 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_351_clock),
    .reset(SaturatingCounter_351_reset),
    .io_enable(SaturatingCounter_351_io_enable),
    .io_value(SaturatingCounter_351_io_value)
  );
  SaturatingCounter SaturatingCounter_352 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_352_clock),
    .reset(SaturatingCounter_352_reset),
    .io_enable(SaturatingCounter_352_io_enable),
    .io_value(SaturatingCounter_352_io_value)
  );
  SaturatingCounter SaturatingCounter_353 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_353_clock),
    .reset(SaturatingCounter_353_reset),
    .io_enable(SaturatingCounter_353_io_enable),
    .io_value(SaturatingCounter_353_io_value)
  );
  SaturatingCounter SaturatingCounter_354 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_354_clock),
    .reset(SaturatingCounter_354_reset),
    .io_enable(SaturatingCounter_354_io_enable),
    .io_value(SaturatingCounter_354_io_value)
  );
  SaturatingCounter SaturatingCounter_355 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_355_clock),
    .reset(SaturatingCounter_355_reset),
    .io_enable(SaturatingCounter_355_io_enable),
    .io_value(SaturatingCounter_355_io_value)
  );
  SaturatingCounter SaturatingCounter_356 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_356_clock),
    .reset(SaturatingCounter_356_reset),
    .io_enable(SaturatingCounter_356_io_enable),
    .io_value(SaturatingCounter_356_io_value)
  );
  SaturatingCounter SaturatingCounter_357 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_357_clock),
    .reset(SaturatingCounter_357_reset),
    .io_enable(SaturatingCounter_357_io_enable),
    .io_value(SaturatingCounter_357_io_value)
  );
  SaturatingCounter SaturatingCounter_358 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_358_clock),
    .reset(SaturatingCounter_358_reset),
    .io_enable(SaturatingCounter_358_io_enable),
    .io_value(SaturatingCounter_358_io_value)
  );
  SaturatingCounter SaturatingCounter_359 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_359_clock),
    .reset(SaturatingCounter_359_reset),
    .io_enable(SaturatingCounter_359_io_enable),
    .io_value(SaturatingCounter_359_io_value)
  );
  SaturatingCounter SaturatingCounter_360 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_360_clock),
    .reset(SaturatingCounter_360_reset),
    .io_enable(SaturatingCounter_360_io_enable),
    .io_value(SaturatingCounter_360_io_value)
  );
  SaturatingCounter SaturatingCounter_361 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_361_clock),
    .reset(SaturatingCounter_361_reset),
    .io_enable(SaturatingCounter_361_io_enable),
    .io_value(SaturatingCounter_361_io_value)
  );
  SaturatingCounter SaturatingCounter_362 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_362_clock),
    .reset(SaturatingCounter_362_reset),
    .io_enable(SaturatingCounter_362_io_enable),
    .io_value(SaturatingCounter_362_io_value)
  );
  SaturatingCounter SaturatingCounter_363 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_363_clock),
    .reset(SaturatingCounter_363_reset),
    .io_enable(SaturatingCounter_363_io_enable),
    .io_value(SaturatingCounter_363_io_value)
  );
  SaturatingCounter SaturatingCounter_364 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_364_clock),
    .reset(SaturatingCounter_364_reset),
    .io_enable(SaturatingCounter_364_io_enable),
    .io_value(SaturatingCounter_364_io_value)
  );
  SaturatingCounter SaturatingCounter_365 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_365_clock),
    .reset(SaturatingCounter_365_reset),
    .io_enable(SaturatingCounter_365_io_enable),
    .io_value(SaturatingCounter_365_io_value)
  );
  SaturatingCounter SaturatingCounter_366 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_366_clock),
    .reset(SaturatingCounter_366_reset),
    .io_enable(SaturatingCounter_366_io_enable),
    .io_value(SaturatingCounter_366_io_value)
  );
  SaturatingCounter SaturatingCounter_367 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_367_clock),
    .reset(SaturatingCounter_367_reset),
    .io_enable(SaturatingCounter_367_io_enable),
    .io_value(SaturatingCounter_367_io_value)
  );
  SaturatingCounter SaturatingCounter_368 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_368_clock),
    .reset(SaturatingCounter_368_reset),
    .io_enable(SaturatingCounter_368_io_enable),
    .io_value(SaturatingCounter_368_io_value)
  );
  SaturatingCounter SaturatingCounter_369 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_369_clock),
    .reset(SaturatingCounter_369_reset),
    .io_enable(SaturatingCounter_369_io_enable),
    .io_value(SaturatingCounter_369_io_value)
  );
  SaturatingCounter SaturatingCounter_370 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_370_clock),
    .reset(SaturatingCounter_370_reset),
    .io_enable(SaturatingCounter_370_io_enable),
    .io_value(SaturatingCounter_370_io_value)
  );
  SaturatingCounter SaturatingCounter_371 ( // @[coverage.scala 105:33]
    .clock(SaturatingCounter_371_clock),
    .reset(SaturatingCounter_371_reset),
    .io_enable(SaturatingCounter_371_io_enable),
    .io_value(SaturatingCounter_371_io_value)
  );
  SaturatingCounter SaturatingCounter_372 ( // @[coverage.scala 107:33]
    .clock(SaturatingCounter_372_clock),
    .reset(SaturatingCounter_372_reset),
    .io_enable(SaturatingCounter_372_io_enable),
    .io_value(SaturatingCounter_372_io_value)
  );
  assign io_coverage_bytes_0 = {7'h0,SaturatingCounter_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_1 = {_T_12,SaturatingCounter_2_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_2 = {_T_16,SaturatingCounter_4_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_3 = {_T_20,SaturatingCounter_6_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_4 = {_T_24,SaturatingCounter_8_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_5 = {_T_28,SaturatingCounter_10_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_6 = {_T_32,SaturatingCounter_12_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_7 = {_T_36,SaturatingCounter_14_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_8 = {_T_40,SaturatingCounter_16_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_9 = {_T_44,SaturatingCounter_18_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_10 = {_T_48,SaturatingCounter_20_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_11 = {_T_52,SaturatingCounter_22_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_12 = {_T_56,SaturatingCounter_24_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_13 = {_T_60,SaturatingCounter_26_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_14 = {_T_64,SaturatingCounter_28_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_15 = {_T_68,SaturatingCounter_30_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_16 = {_T_72,SaturatingCounter_32_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_17 = {_T_76,SaturatingCounter_34_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_18 = {_T_80,SaturatingCounter_36_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_19 = {_T_84,SaturatingCounter_38_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_20 = {_T_88,SaturatingCounter_40_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_21 = {_T_92,SaturatingCounter_42_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_22 = {_T_96,SaturatingCounter_44_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_23 = {_T_100,SaturatingCounter_46_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_24 = {_T_104,SaturatingCounter_48_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_25 = {_T_108,SaturatingCounter_50_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_26 = {_T_112,SaturatingCounter_52_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_27 = {_T_116,SaturatingCounter_54_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_28 = {_T_120,SaturatingCounter_56_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_29 = {_T_124,SaturatingCounter_58_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_30 = {_T_128,SaturatingCounter_60_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_31 = {_T_132,SaturatingCounter_62_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_32 = {_T_136,SaturatingCounter_64_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_33 = {_T_140,SaturatingCounter_66_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_34 = {_T_144,SaturatingCounter_68_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_35 = {_T_148,SaturatingCounter_70_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_36 = {_T_152,SaturatingCounter_72_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_37 = {_T_156,SaturatingCounter_74_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_38 = {_T_160,SaturatingCounter_76_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_39 = {_T_164,SaturatingCounter_78_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_40 = {_T_168,SaturatingCounter_80_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_41 = {_T_172,SaturatingCounter_82_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_42 = {_T_176,SaturatingCounter_84_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_43 = {_T_180,SaturatingCounter_86_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_44 = {_T_184,SaturatingCounter_88_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_45 = {_T_188,SaturatingCounter_90_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_46 = {_T_192,SaturatingCounter_92_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_47 = {_T_196,SaturatingCounter_94_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_48 = {_T_200,SaturatingCounter_96_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_49 = {_T_204,SaturatingCounter_98_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_50 = {_T_208,SaturatingCounter_100_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_51 = {_T_212,SaturatingCounter_102_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_52 = {_T_216,SaturatingCounter_104_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_53 = {_T_220,SaturatingCounter_106_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_54 = {_T_224,SaturatingCounter_108_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_55 = {_T_228,SaturatingCounter_110_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_56 = {_T_232,SaturatingCounter_112_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_57 = {_T_236,SaturatingCounter_114_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_58 = {_T_240,SaturatingCounter_116_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_59 = {_T_244,SaturatingCounter_118_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_60 = {_T_248,SaturatingCounter_120_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_61 = {_T_252,SaturatingCounter_122_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_62 = {_T_256,SaturatingCounter_124_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_63 = {_T_260,SaturatingCounter_126_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_64 = {_T_264,SaturatingCounter_128_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_65 = {_T_268,SaturatingCounter_130_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_66 = {_T_272,SaturatingCounter_132_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_67 = {_T_276,SaturatingCounter_134_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_68 = {_T_280,SaturatingCounter_136_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_69 = {_T_284,SaturatingCounter_138_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_70 = {_T_288,SaturatingCounter_140_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_71 = {_T_292,SaturatingCounter_142_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_72 = {_T_296,SaturatingCounter_144_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_73 = {_T_300,SaturatingCounter_146_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_74 = {_T_304,SaturatingCounter_148_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_75 = {_T_308,SaturatingCounter_150_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_76 = {_T_312,SaturatingCounter_152_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_77 = {_T_316,SaturatingCounter_154_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_78 = {_T_320,SaturatingCounter_156_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_79 = {_T_324,SaturatingCounter_158_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_80 = {_T_328,SaturatingCounter_160_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_81 = {_T_332,SaturatingCounter_162_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_82 = {_T_336,SaturatingCounter_164_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_83 = {_T_340,SaturatingCounter_166_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_84 = {_T_344,SaturatingCounter_168_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_85 = {_T_348,SaturatingCounter_170_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_86 = {_T_352,SaturatingCounter_172_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_87 = {_T_356,SaturatingCounter_174_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_88 = {_T_360,SaturatingCounter_176_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_89 = {_T_364,SaturatingCounter_178_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_90 = {_T_368,SaturatingCounter_180_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_91 = {_T_372,SaturatingCounter_182_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_92 = {_T_376,SaturatingCounter_184_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_93 = {_T_380,SaturatingCounter_186_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_94 = {_T_384,SaturatingCounter_188_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_95 = {_T_388,SaturatingCounter_190_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_96 = {_T_392,SaturatingCounter_192_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_97 = {_T_396,SaturatingCounter_194_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_98 = {_T_400,SaturatingCounter_196_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_99 = {_T_404,SaturatingCounter_198_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_100 = {_T_408,SaturatingCounter_200_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_101 = {_T_412,SaturatingCounter_202_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_102 = {_T_416,SaturatingCounter_204_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_103 = {_T_420,SaturatingCounter_206_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_104 = {_T_424,SaturatingCounter_208_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_105 = {_T_428,SaturatingCounter_210_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_106 = {_T_432,SaturatingCounter_212_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_107 = {_T_436,SaturatingCounter_214_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_108 = {_T_440,SaturatingCounter_216_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_109 = {_T_444,SaturatingCounter_218_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_110 = {_T_448,SaturatingCounter_220_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_111 = {_T_452,SaturatingCounter_222_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_112 = {_T_456,SaturatingCounter_224_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_113 = {_T_460,SaturatingCounter_226_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_114 = {_T_464,SaturatingCounter_228_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_115 = {_T_468,SaturatingCounter_230_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_116 = {_T_472,SaturatingCounter_232_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_117 = {_T_476,SaturatingCounter_234_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_118 = {_T_480,SaturatingCounter_236_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_119 = {_T_484,SaturatingCounter_238_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_120 = {_T_488,SaturatingCounter_240_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_121 = {_T_492,SaturatingCounter_242_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_122 = {_T_496,SaturatingCounter_244_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_123 = {_T_500,SaturatingCounter_246_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_124 = {_T_504,SaturatingCounter_248_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_125 = {_T_508,SaturatingCounter_250_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_126 = {_T_512,SaturatingCounter_252_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_127 = {_T_516,SaturatingCounter_254_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_128 = {_T_520,SaturatingCounter_256_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_129 = {_T_524,SaturatingCounter_258_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_130 = {_T_528,SaturatingCounter_260_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_131 = {_T_532,SaturatingCounter_262_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_132 = {_T_536,SaturatingCounter_264_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_133 = {_T_540,SaturatingCounter_266_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_134 = {_T_544,SaturatingCounter_268_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_135 = {_T_548,SaturatingCounter_270_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_136 = {_T_552,SaturatingCounter_272_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_137 = {_T_556,SaturatingCounter_274_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_138 = {_T_560,SaturatingCounter_276_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_139 = {_T_564,SaturatingCounter_278_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_140 = {_T_568,SaturatingCounter_280_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_141 = {_T_572,SaturatingCounter_282_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_142 = {_T_576,SaturatingCounter_284_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_143 = {_T_580,SaturatingCounter_286_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_144 = {_T_584,SaturatingCounter_288_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_145 = {_T_588,SaturatingCounter_290_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_146 = {_T_592,SaturatingCounter_292_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_147 = {_T_596,SaturatingCounter_294_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_148 = {_T_600,SaturatingCounter_296_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_149 = {_T_604,SaturatingCounter_298_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_150 = {_T_608,SaturatingCounter_300_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_151 = {_T_612,SaturatingCounter_302_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_152 = {_T_616,SaturatingCounter_304_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_153 = {_T_620,SaturatingCounter_306_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_154 = {_T_624,SaturatingCounter_308_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_155 = {_T_628,SaturatingCounter_310_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_156 = {_T_632,SaturatingCounter_312_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_157 = {_T_636,SaturatingCounter_314_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_158 = {_T_640,SaturatingCounter_316_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_159 = {_T_644,SaturatingCounter_318_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_160 = {_T_648,SaturatingCounter_320_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_161 = {_T_652,SaturatingCounter_322_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_162 = {_T_656,SaturatingCounter_324_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_163 = {_T_660,SaturatingCounter_326_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_164 = {_T_664,SaturatingCounter_328_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_165 = {_T_668,SaturatingCounter_330_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_166 = {_T_672,SaturatingCounter_332_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_167 = {_T_676,SaturatingCounter_334_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_168 = {_T_680,SaturatingCounter_336_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_169 = {_T_684,SaturatingCounter_338_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_170 = {_T_688,SaturatingCounter_340_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_171 = {_T_692,SaturatingCounter_342_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_172 = {_T_696,SaturatingCounter_344_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_173 = {_T_700,SaturatingCounter_346_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_174 = {_T_704,SaturatingCounter_348_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_175 = {_T_708,SaturatingCounter_350_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_176 = {_T_712,SaturatingCounter_352_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_177 = {_T_716,SaturatingCounter_354_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_178 = {_T_720,SaturatingCounter_356_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_179 = {_T_724,SaturatingCounter_358_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_180 = {_T_728,SaturatingCounter_360_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_181 = {_T_732,SaturatingCounter_362_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_182 = {_T_736,SaturatingCounter_364_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_183 = {_T_740,SaturatingCounter_366_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_184 = {_T_744,SaturatingCounter_368_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_185 = {_T_748,SaturatingCounter_370_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_186 = {_T_752,SaturatingCounter_372_io_value}; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_187 = 8'h0; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_188 = 8'h0; // @[VerilatorHarness.scala 66:27]
  assign io_coverage_bytes_189 = 8'h0; // @[VerilatorHarness.scala 66:27]
  assign dut_clock = clock;
  assign dut_reset = reset;
  assign dut_io_meta_reset = io_meta_reset; // @[VerilatorHarness.scala 43:27]
  assign dut_io_inputs = input_bytes[63:29]; // @[VerilatorHarness.scala 48:23]
  assign SaturatingCounter_clock = clock;
  assign SaturatingCounter_reset = reset;
  assign SaturatingCounter_io_enable = dut_io_coverage_0; // @[coverage.scala 122:33]
  assign SaturatingCounter_1_clock = clock;
  assign SaturatingCounter_1_reset = reset;
  assign SaturatingCounter_1_io_enable = dut_io_coverage_1; // @[coverage.scala 106:31]
  assign SaturatingCounter_2_clock = clock;
  assign SaturatingCounter_2_reset = reset;
  assign SaturatingCounter_2_io_enable = ~dut_io_coverage_1; // @[coverage.scala 108:31]
  assign SaturatingCounter_3_clock = clock;
  assign SaturatingCounter_3_reset = reset;
  assign SaturatingCounter_3_io_enable = dut_io_coverage_2; // @[coverage.scala 106:31]
  assign SaturatingCounter_4_clock = clock;
  assign SaturatingCounter_4_reset = reset;
  assign SaturatingCounter_4_io_enable = ~dut_io_coverage_2; // @[coverage.scala 108:31]
  assign SaturatingCounter_5_clock = clock;
  assign SaturatingCounter_5_reset = reset;
  assign SaturatingCounter_5_io_enable = dut_io_coverage_3; // @[coverage.scala 106:31]
  assign SaturatingCounter_6_clock = clock;
  assign SaturatingCounter_6_reset = reset;
  assign SaturatingCounter_6_io_enable = ~dut_io_coverage_3; // @[coverage.scala 108:31]
  assign SaturatingCounter_7_clock = clock;
  assign SaturatingCounter_7_reset = reset;
  assign SaturatingCounter_7_io_enable = dut_io_coverage_4; // @[coverage.scala 106:31]
  assign SaturatingCounter_8_clock = clock;
  assign SaturatingCounter_8_reset = reset;
  assign SaturatingCounter_8_io_enable = ~dut_io_coverage_4; // @[coverage.scala 108:31]
  assign SaturatingCounter_9_clock = clock;
  assign SaturatingCounter_9_reset = reset;
  assign SaturatingCounter_9_io_enable = dut_io_coverage_5; // @[coverage.scala 106:31]
  assign SaturatingCounter_10_clock = clock;
  assign SaturatingCounter_10_reset = reset;
  assign SaturatingCounter_10_io_enable = ~dut_io_coverage_5; // @[coverage.scala 108:31]
  assign SaturatingCounter_11_clock = clock;
  assign SaturatingCounter_11_reset = reset;
  assign SaturatingCounter_11_io_enable = dut_io_coverage_6; // @[coverage.scala 106:31]
  assign SaturatingCounter_12_clock = clock;
  assign SaturatingCounter_12_reset = reset;
  assign SaturatingCounter_12_io_enable = ~dut_io_coverage_6; // @[coverage.scala 108:31]
  assign SaturatingCounter_13_clock = clock;
  assign SaturatingCounter_13_reset = reset;
  assign SaturatingCounter_13_io_enable = dut_io_coverage_7; // @[coverage.scala 106:31]
  assign SaturatingCounter_14_clock = clock;
  assign SaturatingCounter_14_reset = reset;
  assign SaturatingCounter_14_io_enable = ~dut_io_coverage_7; // @[coverage.scala 108:31]
  assign SaturatingCounter_15_clock = clock;
  assign SaturatingCounter_15_reset = reset;
  assign SaturatingCounter_15_io_enable = dut_io_coverage_8; // @[coverage.scala 106:31]
  assign SaturatingCounter_16_clock = clock;
  assign SaturatingCounter_16_reset = reset;
  assign SaturatingCounter_16_io_enable = ~dut_io_coverage_8; // @[coverage.scala 108:31]
  assign SaturatingCounter_17_clock = clock;
  assign SaturatingCounter_17_reset = reset;
  assign SaturatingCounter_17_io_enable = dut_io_coverage_9; // @[coverage.scala 106:31]
  assign SaturatingCounter_18_clock = clock;
  assign SaturatingCounter_18_reset = reset;
  assign SaturatingCounter_18_io_enable = ~dut_io_coverage_9; // @[coverage.scala 108:31]
  assign SaturatingCounter_19_clock = clock;
  assign SaturatingCounter_19_reset = reset;
  assign SaturatingCounter_19_io_enable = dut_io_coverage_10; // @[coverage.scala 106:31]
  assign SaturatingCounter_20_clock = clock;
  assign SaturatingCounter_20_reset = reset;
  assign SaturatingCounter_20_io_enable = ~dut_io_coverage_10; // @[coverage.scala 108:31]
  assign SaturatingCounter_21_clock = clock;
  assign SaturatingCounter_21_reset = reset;
  assign SaturatingCounter_21_io_enable = dut_io_coverage_11; // @[coverage.scala 106:31]
  assign SaturatingCounter_22_clock = clock;
  assign SaturatingCounter_22_reset = reset;
  assign SaturatingCounter_22_io_enable = ~dut_io_coverage_11; // @[coverage.scala 108:31]
  assign SaturatingCounter_23_clock = clock;
  assign SaturatingCounter_23_reset = reset;
  assign SaturatingCounter_23_io_enable = dut_io_coverage_12; // @[coverage.scala 106:31]
  assign SaturatingCounter_24_clock = clock;
  assign SaturatingCounter_24_reset = reset;
  assign SaturatingCounter_24_io_enable = ~dut_io_coverage_12; // @[coverage.scala 108:31]
  assign SaturatingCounter_25_clock = clock;
  assign SaturatingCounter_25_reset = reset;
  assign SaturatingCounter_25_io_enable = dut_io_coverage_13; // @[coverage.scala 106:31]
  assign SaturatingCounter_26_clock = clock;
  assign SaturatingCounter_26_reset = reset;
  assign SaturatingCounter_26_io_enable = ~dut_io_coverage_13; // @[coverage.scala 108:31]
  assign SaturatingCounter_27_clock = clock;
  assign SaturatingCounter_27_reset = reset;
  assign SaturatingCounter_27_io_enable = dut_io_coverage_14; // @[coverage.scala 106:31]
  assign SaturatingCounter_28_clock = clock;
  assign SaturatingCounter_28_reset = reset;
  assign SaturatingCounter_28_io_enable = ~dut_io_coverage_14; // @[coverage.scala 108:31]
  assign SaturatingCounter_29_clock = clock;
  assign SaturatingCounter_29_reset = reset;
  assign SaturatingCounter_29_io_enable = dut_io_coverage_15; // @[coverage.scala 106:31]
  assign SaturatingCounter_30_clock = clock;
  assign SaturatingCounter_30_reset = reset;
  assign SaturatingCounter_30_io_enable = ~dut_io_coverage_15; // @[coverage.scala 108:31]
  assign SaturatingCounter_31_clock = clock;
  assign SaturatingCounter_31_reset = reset;
  assign SaturatingCounter_31_io_enable = dut_io_coverage_16; // @[coverage.scala 106:31]
  assign SaturatingCounter_32_clock = clock;
  assign SaturatingCounter_32_reset = reset;
  assign SaturatingCounter_32_io_enable = ~dut_io_coverage_16; // @[coverage.scala 108:31]
  assign SaturatingCounter_33_clock = clock;
  assign SaturatingCounter_33_reset = reset;
  assign SaturatingCounter_33_io_enable = dut_io_coverage_17; // @[coverage.scala 106:31]
  assign SaturatingCounter_34_clock = clock;
  assign SaturatingCounter_34_reset = reset;
  assign SaturatingCounter_34_io_enable = ~dut_io_coverage_17; // @[coverage.scala 108:31]
  assign SaturatingCounter_35_clock = clock;
  assign SaturatingCounter_35_reset = reset;
  assign SaturatingCounter_35_io_enable = dut_io_coverage_18; // @[coverage.scala 106:31]
  assign SaturatingCounter_36_clock = clock;
  assign SaturatingCounter_36_reset = reset;
  assign SaturatingCounter_36_io_enable = ~dut_io_coverage_18; // @[coverage.scala 108:31]
  assign SaturatingCounter_37_clock = clock;
  assign SaturatingCounter_37_reset = reset;
  assign SaturatingCounter_37_io_enable = dut_io_coverage_19; // @[coverage.scala 106:31]
  assign SaturatingCounter_38_clock = clock;
  assign SaturatingCounter_38_reset = reset;
  assign SaturatingCounter_38_io_enable = ~dut_io_coverage_19; // @[coverage.scala 108:31]
  assign SaturatingCounter_39_clock = clock;
  assign SaturatingCounter_39_reset = reset;
  assign SaturatingCounter_39_io_enable = dut_io_coverage_20; // @[coverage.scala 106:31]
  assign SaturatingCounter_40_clock = clock;
  assign SaturatingCounter_40_reset = reset;
  assign SaturatingCounter_40_io_enable = ~dut_io_coverage_20; // @[coverage.scala 108:31]
  assign SaturatingCounter_41_clock = clock;
  assign SaturatingCounter_41_reset = reset;
  assign SaturatingCounter_41_io_enable = dut_io_coverage_21; // @[coverage.scala 106:31]
  assign SaturatingCounter_42_clock = clock;
  assign SaturatingCounter_42_reset = reset;
  assign SaturatingCounter_42_io_enable = ~dut_io_coverage_21; // @[coverage.scala 108:31]
  assign SaturatingCounter_43_clock = clock;
  assign SaturatingCounter_43_reset = reset;
  assign SaturatingCounter_43_io_enable = dut_io_coverage_22; // @[coverage.scala 106:31]
  assign SaturatingCounter_44_clock = clock;
  assign SaturatingCounter_44_reset = reset;
  assign SaturatingCounter_44_io_enable = ~dut_io_coverage_22; // @[coverage.scala 108:31]
  assign SaturatingCounter_45_clock = clock;
  assign SaturatingCounter_45_reset = reset;
  assign SaturatingCounter_45_io_enable = dut_io_coverage_23; // @[coverage.scala 106:31]
  assign SaturatingCounter_46_clock = clock;
  assign SaturatingCounter_46_reset = reset;
  assign SaturatingCounter_46_io_enable = ~dut_io_coverage_23; // @[coverage.scala 108:31]
  assign SaturatingCounter_47_clock = clock;
  assign SaturatingCounter_47_reset = reset;
  assign SaturatingCounter_47_io_enable = dut_io_coverage_24; // @[coverage.scala 106:31]
  assign SaturatingCounter_48_clock = clock;
  assign SaturatingCounter_48_reset = reset;
  assign SaturatingCounter_48_io_enable = ~dut_io_coverage_24; // @[coverage.scala 108:31]
  assign SaturatingCounter_49_clock = clock;
  assign SaturatingCounter_49_reset = reset;
  assign SaturatingCounter_49_io_enable = dut_io_coverage_25; // @[coverage.scala 106:31]
  assign SaturatingCounter_50_clock = clock;
  assign SaturatingCounter_50_reset = reset;
  assign SaturatingCounter_50_io_enable = ~dut_io_coverage_25; // @[coverage.scala 108:31]
  assign SaturatingCounter_51_clock = clock;
  assign SaturatingCounter_51_reset = reset;
  assign SaturatingCounter_51_io_enable = dut_io_coverage_26; // @[coverage.scala 106:31]
  assign SaturatingCounter_52_clock = clock;
  assign SaturatingCounter_52_reset = reset;
  assign SaturatingCounter_52_io_enable = ~dut_io_coverage_26; // @[coverage.scala 108:31]
  assign SaturatingCounter_53_clock = clock;
  assign SaturatingCounter_53_reset = reset;
  assign SaturatingCounter_53_io_enable = dut_io_coverage_27; // @[coverage.scala 106:31]
  assign SaturatingCounter_54_clock = clock;
  assign SaturatingCounter_54_reset = reset;
  assign SaturatingCounter_54_io_enable = ~dut_io_coverage_27; // @[coverage.scala 108:31]
  assign SaturatingCounter_55_clock = clock;
  assign SaturatingCounter_55_reset = reset;
  assign SaturatingCounter_55_io_enable = dut_io_coverage_28; // @[coverage.scala 106:31]
  assign SaturatingCounter_56_clock = clock;
  assign SaturatingCounter_56_reset = reset;
  assign SaturatingCounter_56_io_enable = ~dut_io_coverage_28; // @[coverage.scala 108:31]
  assign SaturatingCounter_57_clock = clock;
  assign SaturatingCounter_57_reset = reset;
  assign SaturatingCounter_57_io_enable = dut_io_coverage_29; // @[coverage.scala 106:31]
  assign SaturatingCounter_58_clock = clock;
  assign SaturatingCounter_58_reset = reset;
  assign SaturatingCounter_58_io_enable = ~dut_io_coverage_29; // @[coverage.scala 108:31]
  assign SaturatingCounter_59_clock = clock;
  assign SaturatingCounter_59_reset = reset;
  assign SaturatingCounter_59_io_enable = dut_io_coverage_30; // @[coverage.scala 106:31]
  assign SaturatingCounter_60_clock = clock;
  assign SaturatingCounter_60_reset = reset;
  assign SaturatingCounter_60_io_enable = ~dut_io_coverage_30; // @[coverage.scala 108:31]
  assign SaturatingCounter_61_clock = clock;
  assign SaturatingCounter_61_reset = reset;
  assign SaturatingCounter_61_io_enable = dut_io_coverage_31; // @[coverage.scala 106:31]
  assign SaturatingCounter_62_clock = clock;
  assign SaturatingCounter_62_reset = reset;
  assign SaturatingCounter_62_io_enable = ~dut_io_coverage_31; // @[coverage.scala 108:31]
  assign SaturatingCounter_63_clock = clock;
  assign SaturatingCounter_63_reset = reset;
  assign SaturatingCounter_63_io_enable = dut_io_coverage_32; // @[coverage.scala 106:31]
  assign SaturatingCounter_64_clock = clock;
  assign SaturatingCounter_64_reset = reset;
  assign SaturatingCounter_64_io_enable = ~dut_io_coverage_32; // @[coverage.scala 108:31]
  assign SaturatingCounter_65_clock = clock;
  assign SaturatingCounter_65_reset = reset;
  assign SaturatingCounter_65_io_enable = dut_io_coverage_33; // @[coverage.scala 106:31]
  assign SaturatingCounter_66_clock = clock;
  assign SaturatingCounter_66_reset = reset;
  assign SaturatingCounter_66_io_enable = ~dut_io_coverage_33; // @[coverage.scala 108:31]
  assign SaturatingCounter_67_clock = clock;
  assign SaturatingCounter_67_reset = reset;
  assign SaturatingCounter_67_io_enable = dut_io_coverage_34; // @[coverage.scala 106:31]
  assign SaturatingCounter_68_clock = clock;
  assign SaturatingCounter_68_reset = reset;
  assign SaturatingCounter_68_io_enable = ~dut_io_coverage_34; // @[coverage.scala 108:31]
  assign SaturatingCounter_69_clock = clock;
  assign SaturatingCounter_69_reset = reset;
  assign SaturatingCounter_69_io_enable = dut_io_coverage_35; // @[coverage.scala 106:31]
  assign SaturatingCounter_70_clock = clock;
  assign SaturatingCounter_70_reset = reset;
  assign SaturatingCounter_70_io_enable = ~dut_io_coverage_35; // @[coverage.scala 108:31]
  assign SaturatingCounter_71_clock = clock;
  assign SaturatingCounter_71_reset = reset;
  assign SaturatingCounter_71_io_enable = dut_io_coverage_36; // @[coverage.scala 106:31]
  assign SaturatingCounter_72_clock = clock;
  assign SaturatingCounter_72_reset = reset;
  assign SaturatingCounter_72_io_enable = ~dut_io_coverage_36; // @[coverage.scala 108:31]
  assign SaturatingCounter_73_clock = clock;
  assign SaturatingCounter_73_reset = reset;
  assign SaturatingCounter_73_io_enable = dut_io_coverage_37; // @[coverage.scala 106:31]
  assign SaturatingCounter_74_clock = clock;
  assign SaturatingCounter_74_reset = reset;
  assign SaturatingCounter_74_io_enable = ~dut_io_coverage_37; // @[coverage.scala 108:31]
  assign SaturatingCounter_75_clock = clock;
  assign SaturatingCounter_75_reset = reset;
  assign SaturatingCounter_75_io_enable = dut_io_coverage_38; // @[coverage.scala 106:31]
  assign SaturatingCounter_76_clock = clock;
  assign SaturatingCounter_76_reset = reset;
  assign SaturatingCounter_76_io_enable = ~dut_io_coverage_38; // @[coverage.scala 108:31]
  assign SaturatingCounter_77_clock = clock;
  assign SaturatingCounter_77_reset = reset;
  assign SaturatingCounter_77_io_enable = dut_io_coverage_39; // @[coverage.scala 106:31]
  assign SaturatingCounter_78_clock = clock;
  assign SaturatingCounter_78_reset = reset;
  assign SaturatingCounter_78_io_enable = ~dut_io_coverage_39; // @[coverage.scala 108:31]
  assign SaturatingCounter_79_clock = clock;
  assign SaturatingCounter_79_reset = reset;
  assign SaturatingCounter_79_io_enable = dut_io_coverage_40; // @[coverage.scala 106:31]
  assign SaturatingCounter_80_clock = clock;
  assign SaturatingCounter_80_reset = reset;
  assign SaturatingCounter_80_io_enable = ~dut_io_coverage_40; // @[coverage.scala 108:31]
  assign SaturatingCounter_81_clock = clock;
  assign SaturatingCounter_81_reset = reset;
  assign SaturatingCounter_81_io_enable = dut_io_coverage_41; // @[coverage.scala 106:31]
  assign SaturatingCounter_82_clock = clock;
  assign SaturatingCounter_82_reset = reset;
  assign SaturatingCounter_82_io_enable = ~dut_io_coverage_41; // @[coverage.scala 108:31]
  assign SaturatingCounter_83_clock = clock;
  assign SaturatingCounter_83_reset = reset;
  assign SaturatingCounter_83_io_enable = dut_io_coverage_42; // @[coverage.scala 106:31]
  assign SaturatingCounter_84_clock = clock;
  assign SaturatingCounter_84_reset = reset;
  assign SaturatingCounter_84_io_enable = ~dut_io_coverage_42; // @[coverage.scala 108:31]
  assign SaturatingCounter_85_clock = clock;
  assign SaturatingCounter_85_reset = reset;
  assign SaturatingCounter_85_io_enable = dut_io_coverage_43; // @[coverage.scala 106:31]
  assign SaturatingCounter_86_clock = clock;
  assign SaturatingCounter_86_reset = reset;
  assign SaturatingCounter_86_io_enable = ~dut_io_coverage_43; // @[coverage.scala 108:31]
  assign SaturatingCounter_87_clock = clock;
  assign SaturatingCounter_87_reset = reset;
  assign SaturatingCounter_87_io_enable = dut_io_coverage_44; // @[coverage.scala 106:31]
  assign SaturatingCounter_88_clock = clock;
  assign SaturatingCounter_88_reset = reset;
  assign SaturatingCounter_88_io_enable = ~dut_io_coverage_44; // @[coverage.scala 108:31]
  assign SaturatingCounter_89_clock = clock;
  assign SaturatingCounter_89_reset = reset;
  assign SaturatingCounter_89_io_enable = dut_io_coverage_45; // @[coverage.scala 106:31]
  assign SaturatingCounter_90_clock = clock;
  assign SaturatingCounter_90_reset = reset;
  assign SaturatingCounter_90_io_enable = ~dut_io_coverage_45; // @[coverage.scala 108:31]
  assign SaturatingCounter_91_clock = clock;
  assign SaturatingCounter_91_reset = reset;
  assign SaturatingCounter_91_io_enable = dut_io_coverage_46; // @[coverage.scala 106:31]
  assign SaturatingCounter_92_clock = clock;
  assign SaturatingCounter_92_reset = reset;
  assign SaturatingCounter_92_io_enable = ~dut_io_coverage_46; // @[coverage.scala 108:31]
  assign SaturatingCounter_93_clock = clock;
  assign SaturatingCounter_93_reset = reset;
  assign SaturatingCounter_93_io_enable = dut_io_coverage_47; // @[coverage.scala 106:31]
  assign SaturatingCounter_94_clock = clock;
  assign SaturatingCounter_94_reset = reset;
  assign SaturatingCounter_94_io_enable = ~dut_io_coverage_47; // @[coverage.scala 108:31]
  assign SaturatingCounter_95_clock = clock;
  assign SaturatingCounter_95_reset = reset;
  assign SaturatingCounter_95_io_enable = dut_io_coverage_48; // @[coverage.scala 106:31]
  assign SaturatingCounter_96_clock = clock;
  assign SaturatingCounter_96_reset = reset;
  assign SaturatingCounter_96_io_enable = ~dut_io_coverage_48; // @[coverage.scala 108:31]
  assign SaturatingCounter_97_clock = clock;
  assign SaturatingCounter_97_reset = reset;
  assign SaturatingCounter_97_io_enable = dut_io_coverage_49; // @[coverage.scala 106:31]
  assign SaturatingCounter_98_clock = clock;
  assign SaturatingCounter_98_reset = reset;
  assign SaturatingCounter_98_io_enable = ~dut_io_coverage_49; // @[coverage.scala 108:31]
  assign SaturatingCounter_99_clock = clock;
  assign SaturatingCounter_99_reset = reset;
  assign SaturatingCounter_99_io_enable = dut_io_coverage_50; // @[coverage.scala 106:31]
  assign SaturatingCounter_100_clock = clock;
  assign SaturatingCounter_100_reset = reset;
  assign SaturatingCounter_100_io_enable = ~dut_io_coverage_50; // @[coverage.scala 108:31]
  assign SaturatingCounter_101_clock = clock;
  assign SaturatingCounter_101_reset = reset;
  assign SaturatingCounter_101_io_enable = dut_io_coverage_51; // @[coverage.scala 106:31]
  assign SaturatingCounter_102_clock = clock;
  assign SaturatingCounter_102_reset = reset;
  assign SaturatingCounter_102_io_enable = ~dut_io_coverage_51; // @[coverage.scala 108:31]
  assign SaturatingCounter_103_clock = clock;
  assign SaturatingCounter_103_reset = reset;
  assign SaturatingCounter_103_io_enable = dut_io_coverage_52; // @[coverage.scala 106:31]
  assign SaturatingCounter_104_clock = clock;
  assign SaturatingCounter_104_reset = reset;
  assign SaturatingCounter_104_io_enable = ~dut_io_coverage_52; // @[coverage.scala 108:31]
  assign SaturatingCounter_105_clock = clock;
  assign SaturatingCounter_105_reset = reset;
  assign SaturatingCounter_105_io_enable = dut_io_coverage_53; // @[coverage.scala 106:31]
  assign SaturatingCounter_106_clock = clock;
  assign SaturatingCounter_106_reset = reset;
  assign SaturatingCounter_106_io_enable = ~dut_io_coverage_53; // @[coverage.scala 108:31]
  assign SaturatingCounter_107_clock = clock;
  assign SaturatingCounter_107_reset = reset;
  assign SaturatingCounter_107_io_enable = dut_io_coverage_54; // @[coverage.scala 106:31]
  assign SaturatingCounter_108_clock = clock;
  assign SaturatingCounter_108_reset = reset;
  assign SaturatingCounter_108_io_enable = ~dut_io_coverage_54; // @[coverage.scala 108:31]
  assign SaturatingCounter_109_clock = clock;
  assign SaturatingCounter_109_reset = reset;
  assign SaturatingCounter_109_io_enable = dut_io_coverage_55; // @[coverage.scala 106:31]
  assign SaturatingCounter_110_clock = clock;
  assign SaturatingCounter_110_reset = reset;
  assign SaturatingCounter_110_io_enable = ~dut_io_coverage_55; // @[coverage.scala 108:31]
  assign SaturatingCounter_111_clock = clock;
  assign SaturatingCounter_111_reset = reset;
  assign SaturatingCounter_111_io_enable = dut_io_coverage_56; // @[coverage.scala 106:31]
  assign SaturatingCounter_112_clock = clock;
  assign SaturatingCounter_112_reset = reset;
  assign SaturatingCounter_112_io_enable = ~dut_io_coverage_56; // @[coverage.scala 108:31]
  assign SaturatingCounter_113_clock = clock;
  assign SaturatingCounter_113_reset = reset;
  assign SaturatingCounter_113_io_enable = dut_io_coverage_57; // @[coverage.scala 106:31]
  assign SaturatingCounter_114_clock = clock;
  assign SaturatingCounter_114_reset = reset;
  assign SaturatingCounter_114_io_enable = ~dut_io_coverage_57; // @[coverage.scala 108:31]
  assign SaturatingCounter_115_clock = clock;
  assign SaturatingCounter_115_reset = reset;
  assign SaturatingCounter_115_io_enable = dut_io_coverage_58; // @[coverage.scala 106:31]
  assign SaturatingCounter_116_clock = clock;
  assign SaturatingCounter_116_reset = reset;
  assign SaturatingCounter_116_io_enable = ~dut_io_coverage_58; // @[coverage.scala 108:31]
  assign SaturatingCounter_117_clock = clock;
  assign SaturatingCounter_117_reset = reset;
  assign SaturatingCounter_117_io_enable = dut_io_coverage_59; // @[coverage.scala 106:31]
  assign SaturatingCounter_118_clock = clock;
  assign SaturatingCounter_118_reset = reset;
  assign SaturatingCounter_118_io_enable = ~dut_io_coverage_59; // @[coverage.scala 108:31]
  assign SaturatingCounter_119_clock = clock;
  assign SaturatingCounter_119_reset = reset;
  assign SaturatingCounter_119_io_enable = dut_io_coverage_60; // @[coverage.scala 106:31]
  assign SaturatingCounter_120_clock = clock;
  assign SaturatingCounter_120_reset = reset;
  assign SaturatingCounter_120_io_enable = ~dut_io_coverage_60; // @[coverage.scala 108:31]
  assign SaturatingCounter_121_clock = clock;
  assign SaturatingCounter_121_reset = reset;
  assign SaturatingCounter_121_io_enable = dut_io_coverage_61; // @[coverage.scala 106:31]
  assign SaturatingCounter_122_clock = clock;
  assign SaturatingCounter_122_reset = reset;
  assign SaturatingCounter_122_io_enable = ~dut_io_coverage_61; // @[coverage.scala 108:31]
  assign SaturatingCounter_123_clock = clock;
  assign SaturatingCounter_123_reset = reset;
  assign SaturatingCounter_123_io_enable = dut_io_coverage_62; // @[coverage.scala 106:31]
  assign SaturatingCounter_124_clock = clock;
  assign SaturatingCounter_124_reset = reset;
  assign SaturatingCounter_124_io_enable = ~dut_io_coverage_62; // @[coverage.scala 108:31]
  assign SaturatingCounter_125_clock = clock;
  assign SaturatingCounter_125_reset = reset;
  assign SaturatingCounter_125_io_enable = dut_io_coverage_63; // @[coverage.scala 106:31]
  assign SaturatingCounter_126_clock = clock;
  assign SaturatingCounter_126_reset = reset;
  assign SaturatingCounter_126_io_enable = ~dut_io_coverage_63; // @[coverage.scala 108:31]
  assign SaturatingCounter_127_clock = clock;
  assign SaturatingCounter_127_reset = reset;
  assign SaturatingCounter_127_io_enable = dut_io_coverage_64; // @[coverage.scala 106:31]
  assign SaturatingCounter_128_clock = clock;
  assign SaturatingCounter_128_reset = reset;
  assign SaturatingCounter_128_io_enable = ~dut_io_coverage_64; // @[coverage.scala 108:31]
  assign SaturatingCounter_129_clock = clock;
  assign SaturatingCounter_129_reset = reset;
  assign SaturatingCounter_129_io_enable = dut_io_coverage_65; // @[coverage.scala 106:31]
  assign SaturatingCounter_130_clock = clock;
  assign SaturatingCounter_130_reset = reset;
  assign SaturatingCounter_130_io_enable = ~dut_io_coverage_65; // @[coverage.scala 108:31]
  assign SaturatingCounter_131_clock = clock;
  assign SaturatingCounter_131_reset = reset;
  assign SaturatingCounter_131_io_enable = dut_io_coverage_66; // @[coverage.scala 106:31]
  assign SaturatingCounter_132_clock = clock;
  assign SaturatingCounter_132_reset = reset;
  assign SaturatingCounter_132_io_enable = ~dut_io_coverage_66; // @[coverage.scala 108:31]
  assign SaturatingCounter_133_clock = clock;
  assign SaturatingCounter_133_reset = reset;
  assign SaturatingCounter_133_io_enable = dut_io_coverage_67; // @[coverage.scala 106:31]
  assign SaturatingCounter_134_clock = clock;
  assign SaturatingCounter_134_reset = reset;
  assign SaturatingCounter_134_io_enable = ~dut_io_coverage_67; // @[coverage.scala 108:31]
  assign SaturatingCounter_135_clock = clock;
  assign SaturatingCounter_135_reset = reset;
  assign SaturatingCounter_135_io_enable = dut_io_coverage_68; // @[coverage.scala 106:31]
  assign SaturatingCounter_136_clock = clock;
  assign SaturatingCounter_136_reset = reset;
  assign SaturatingCounter_136_io_enable = ~dut_io_coverage_68; // @[coverage.scala 108:31]
  assign SaturatingCounter_137_clock = clock;
  assign SaturatingCounter_137_reset = reset;
  assign SaturatingCounter_137_io_enable = dut_io_coverage_69; // @[coverage.scala 106:31]
  assign SaturatingCounter_138_clock = clock;
  assign SaturatingCounter_138_reset = reset;
  assign SaturatingCounter_138_io_enable = ~dut_io_coverage_69; // @[coverage.scala 108:31]
  assign SaturatingCounter_139_clock = clock;
  assign SaturatingCounter_139_reset = reset;
  assign SaturatingCounter_139_io_enable = dut_io_coverage_70; // @[coverage.scala 106:31]
  assign SaturatingCounter_140_clock = clock;
  assign SaturatingCounter_140_reset = reset;
  assign SaturatingCounter_140_io_enable = ~dut_io_coverage_70; // @[coverage.scala 108:31]
  assign SaturatingCounter_141_clock = clock;
  assign SaturatingCounter_141_reset = reset;
  assign SaturatingCounter_141_io_enable = dut_io_coverage_71; // @[coverage.scala 106:31]
  assign SaturatingCounter_142_clock = clock;
  assign SaturatingCounter_142_reset = reset;
  assign SaturatingCounter_142_io_enable = ~dut_io_coverage_71; // @[coverage.scala 108:31]
  assign SaturatingCounter_143_clock = clock;
  assign SaturatingCounter_143_reset = reset;
  assign SaturatingCounter_143_io_enable = dut_io_coverage_72; // @[coverage.scala 106:31]
  assign SaturatingCounter_144_clock = clock;
  assign SaturatingCounter_144_reset = reset;
  assign SaturatingCounter_144_io_enable = ~dut_io_coverage_72; // @[coverage.scala 108:31]
  assign SaturatingCounter_145_clock = clock;
  assign SaturatingCounter_145_reset = reset;
  assign SaturatingCounter_145_io_enable = dut_io_coverage_73; // @[coverage.scala 106:31]
  assign SaturatingCounter_146_clock = clock;
  assign SaturatingCounter_146_reset = reset;
  assign SaturatingCounter_146_io_enable = ~dut_io_coverage_73; // @[coverage.scala 108:31]
  assign SaturatingCounter_147_clock = clock;
  assign SaturatingCounter_147_reset = reset;
  assign SaturatingCounter_147_io_enable = dut_io_coverage_74; // @[coverage.scala 106:31]
  assign SaturatingCounter_148_clock = clock;
  assign SaturatingCounter_148_reset = reset;
  assign SaturatingCounter_148_io_enable = ~dut_io_coverage_74; // @[coverage.scala 108:31]
  assign SaturatingCounter_149_clock = clock;
  assign SaturatingCounter_149_reset = reset;
  assign SaturatingCounter_149_io_enable = dut_io_coverage_75; // @[coverage.scala 106:31]
  assign SaturatingCounter_150_clock = clock;
  assign SaturatingCounter_150_reset = reset;
  assign SaturatingCounter_150_io_enable = ~dut_io_coverage_75; // @[coverage.scala 108:31]
  assign SaturatingCounter_151_clock = clock;
  assign SaturatingCounter_151_reset = reset;
  assign SaturatingCounter_151_io_enable = dut_io_coverage_76; // @[coverage.scala 106:31]
  assign SaturatingCounter_152_clock = clock;
  assign SaturatingCounter_152_reset = reset;
  assign SaturatingCounter_152_io_enable = ~dut_io_coverage_76; // @[coverage.scala 108:31]
  assign SaturatingCounter_153_clock = clock;
  assign SaturatingCounter_153_reset = reset;
  assign SaturatingCounter_153_io_enable = dut_io_coverage_77; // @[coverage.scala 106:31]
  assign SaturatingCounter_154_clock = clock;
  assign SaturatingCounter_154_reset = reset;
  assign SaturatingCounter_154_io_enable = ~dut_io_coverage_77; // @[coverage.scala 108:31]
  assign SaturatingCounter_155_clock = clock;
  assign SaturatingCounter_155_reset = reset;
  assign SaturatingCounter_155_io_enable = dut_io_coverage_78; // @[coverage.scala 106:31]
  assign SaturatingCounter_156_clock = clock;
  assign SaturatingCounter_156_reset = reset;
  assign SaturatingCounter_156_io_enable = ~dut_io_coverage_78; // @[coverage.scala 108:31]
  assign SaturatingCounter_157_clock = clock;
  assign SaturatingCounter_157_reset = reset;
  assign SaturatingCounter_157_io_enable = dut_io_coverage_79; // @[coverage.scala 106:31]
  assign SaturatingCounter_158_clock = clock;
  assign SaturatingCounter_158_reset = reset;
  assign SaturatingCounter_158_io_enable = ~dut_io_coverage_79; // @[coverage.scala 108:31]
  assign SaturatingCounter_159_clock = clock;
  assign SaturatingCounter_159_reset = reset;
  assign SaturatingCounter_159_io_enable = dut_io_coverage_80; // @[coverage.scala 106:31]
  assign SaturatingCounter_160_clock = clock;
  assign SaturatingCounter_160_reset = reset;
  assign SaturatingCounter_160_io_enable = ~dut_io_coverage_80; // @[coverage.scala 108:31]
  assign SaturatingCounter_161_clock = clock;
  assign SaturatingCounter_161_reset = reset;
  assign SaturatingCounter_161_io_enable = dut_io_coverage_81; // @[coverage.scala 106:31]
  assign SaturatingCounter_162_clock = clock;
  assign SaturatingCounter_162_reset = reset;
  assign SaturatingCounter_162_io_enable = ~dut_io_coverage_81; // @[coverage.scala 108:31]
  assign SaturatingCounter_163_clock = clock;
  assign SaturatingCounter_163_reset = reset;
  assign SaturatingCounter_163_io_enable = dut_io_coverage_82; // @[coverage.scala 106:31]
  assign SaturatingCounter_164_clock = clock;
  assign SaturatingCounter_164_reset = reset;
  assign SaturatingCounter_164_io_enable = ~dut_io_coverage_82; // @[coverage.scala 108:31]
  assign SaturatingCounter_165_clock = clock;
  assign SaturatingCounter_165_reset = reset;
  assign SaturatingCounter_165_io_enable = dut_io_coverage_83; // @[coverage.scala 106:31]
  assign SaturatingCounter_166_clock = clock;
  assign SaturatingCounter_166_reset = reset;
  assign SaturatingCounter_166_io_enable = ~dut_io_coverage_83; // @[coverage.scala 108:31]
  assign SaturatingCounter_167_clock = clock;
  assign SaturatingCounter_167_reset = reset;
  assign SaturatingCounter_167_io_enable = dut_io_coverage_84; // @[coverage.scala 106:31]
  assign SaturatingCounter_168_clock = clock;
  assign SaturatingCounter_168_reset = reset;
  assign SaturatingCounter_168_io_enable = ~dut_io_coverage_84; // @[coverage.scala 108:31]
  assign SaturatingCounter_169_clock = clock;
  assign SaturatingCounter_169_reset = reset;
  assign SaturatingCounter_169_io_enable = dut_io_coverage_85; // @[coverage.scala 106:31]
  assign SaturatingCounter_170_clock = clock;
  assign SaturatingCounter_170_reset = reset;
  assign SaturatingCounter_170_io_enable = ~dut_io_coverage_85; // @[coverage.scala 108:31]
  assign SaturatingCounter_171_clock = clock;
  assign SaturatingCounter_171_reset = reset;
  assign SaturatingCounter_171_io_enable = dut_io_coverage_86; // @[coverage.scala 106:31]
  assign SaturatingCounter_172_clock = clock;
  assign SaturatingCounter_172_reset = reset;
  assign SaturatingCounter_172_io_enable = ~dut_io_coverage_86; // @[coverage.scala 108:31]
  assign SaturatingCounter_173_clock = clock;
  assign SaturatingCounter_173_reset = reset;
  assign SaturatingCounter_173_io_enable = dut_io_coverage_87; // @[coverage.scala 106:31]
  assign SaturatingCounter_174_clock = clock;
  assign SaturatingCounter_174_reset = reset;
  assign SaturatingCounter_174_io_enable = ~dut_io_coverage_87; // @[coverage.scala 108:31]
  assign SaturatingCounter_175_clock = clock;
  assign SaturatingCounter_175_reset = reset;
  assign SaturatingCounter_175_io_enable = dut_io_coverage_88; // @[coverage.scala 106:31]
  assign SaturatingCounter_176_clock = clock;
  assign SaturatingCounter_176_reset = reset;
  assign SaturatingCounter_176_io_enable = ~dut_io_coverage_88; // @[coverage.scala 108:31]
  assign SaturatingCounter_177_clock = clock;
  assign SaturatingCounter_177_reset = reset;
  assign SaturatingCounter_177_io_enable = dut_io_coverage_89; // @[coverage.scala 106:31]
  assign SaturatingCounter_178_clock = clock;
  assign SaturatingCounter_178_reset = reset;
  assign SaturatingCounter_178_io_enable = ~dut_io_coverage_89; // @[coverage.scala 108:31]
  assign SaturatingCounter_179_clock = clock;
  assign SaturatingCounter_179_reset = reset;
  assign SaturatingCounter_179_io_enable = dut_io_coverage_90; // @[coverage.scala 106:31]
  assign SaturatingCounter_180_clock = clock;
  assign SaturatingCounter_180_reset = reset;
  assign SaturatingCounter_180_io_enable = ~dut_io_coverage_90; // @[coverage.scala 108:31]
  assign SaturatingCounter_181_clock = clock;
  assign SaturatingCounter_181_reset = reset;
  assign SaturatingCounter_181_io_enable = dut_io_coverage_91; // @[coverage.scala 106:31]
  assign SaturatingCounter_182_clock = clock;
  assign SaturatingCounter_182_reset = reset;
  assign SaturatingCounter_182_io_enable = ~dut_io_coverage_91; // @[coverage.scala 108:31]
  assign SaturatingCounter_183_clock = clock;
  assign SaturatingCounter_183_reset = reset;
  assign SaturatingCounter_183_io_enable = dut_io_coverage_92; // @[coverage.scala 106:31]
  assign SaturatingCounter_184_clock = clock;
  assign SaturatingCounter_184_reset = reset;
  assign SaturatingCounter_184_io_enable = ~dut_io_coverage_92; // @[coverage.scala 108:31]
  assign SaturatingCounter_185_clock = clock;
  assign SaturatingCounter_185_reset = reset;
  assign SaturatingCounter_185_io_enable = dut_io_coverage_93; // @[coverage.scala 106:31]
  assign SaturatingCounter_186_clock = clock;
  assign SaturatingCounter_186_reset = reset;
  assign SaturatingCounter_186_io_enable = ~dut_io_coverage_93; // @[coverage.scala 108:31]
  assign SaturatingCounter_187_clock = clock;
  assign SaturatingCounter_187_reset = reset;
  assign SaturatingCounter_187_io_enable = dut_io_coverage_94; // @[coverage.scala 106:31]
  assign SaturatingCounter_188_clock = clock;
  assign SaturatingCounter_188_reset = reset;
  assign SaturatingCounter_188_io_enable = ~dut_io_coverage_94; // @[coverage.scala 108:31]
  assign SaturatingCounter_189_clock = clock;
  assign SaturatingCounter_189_reset = reset;
  assign SaturatingCounter_189_io_enable = dut_io_coverage_95; // @[coverage.scala 106:31]
  assign SaturatingCounter_190_clock = clock;
  assign SaturatingCounter_190_reset = reset;
  assign SaturatingCounter_190_io_enable = ~dut_io_coverage_95; // @[coverage.scala 108:31]
  assign SaturatingCounter_191_clock = clock;
  assign SaturatingCounter_191_reset = reset;
  assign SaturatingCounter_191_io_enable = dut_io_coverage_96; // @[coverage.scala 106:31]
  assign SaturatingCounter_192_clock = clock;
  assign SaturatingCounter_192_reset = reset;
  assign SaturatingCounter_192_io_enable = ~dut_io_coverage_96; // @[coverage.scala 108:31]
  assign SaturatingCounter_193_clock = clock;
  assign SaturatingCounter_193_reset = reset;
  assign SaturatingCounter_193_io_enable = dut_io_coverage_97; // @[coverage.scala 106:31]
  assign SaturatingCounter_194_clock = clock;
  assign SaturatingCounter_194_reset = reset;
  assign SaturatingCounter_194_io_enable = ~dut_io_coverage_97; // @[coverage.scala 108:31]
  assign SaturatingCounter_195_clock = clock;
  assign SaturatingCounter_195_reset = reset;
  assign SaturatingCounter_195_io_enable = dut_io_coverage_98; // @[coverage.scala 106:31]
  assign SaturatingCounter_196_clock = clock;
  assign SaturatingCounter_196_reset = reset;
  assign SaturatingCounter_196_io_enable = ~dut_io_coverage_98; // @[coverage.scala 108:31]
  assign SaturatingCounter_197_clock = clock;
  assign SaturatingCounter_197_reset = reset;
  assign SaturatingCounter_197_io_enable = dut_io_coverage_99; // @[coverage.scala 106:31]
  assign SaturatingCounter_198_clock = clock;
  assign SaturatingCounter_198_reset = reset;
  assign SaturatingCounter_198_io_enable = ~dut_io_coverage_99; // @[coverage.scala 108:31]
  assign SaturatingCounter_199_clock = clock;
  assign SaturatingCounter_199_reset = reset;
  assign SaturatingCounter_199_io_enable = dut_io_coverage_100; // @[coverage.scala 106:31]
  assign SaturatingCounter_200_clock = clock;
  assign SaturatingCounter_200_reset = reset;
  assign SaturatingCounter_200_io_enable = ~dut_io_coverage_100; // @[coverage.scala 108:31]
  assign SaturatingCounter_201_clock = clock;
  assign SaturatingCounter_201_reset = reset;
  assign SaturatingCounter_201_io_enable = dut_io_coverage_101; // @[coverage.scala 106:31]
  assign SaturatingCounter_202_clock = clock;
  assign SaturatingCounter_202_reset = reset;
  assign SaturatingCounter_202_io_enable = ~dut_io_coverage_101; // @[coverage.scala 108:31]
  assign SaturatingCounter_203_clock = clock;
  assign SaturatingCounter_203_reset = reset;
  assign SaturatingCounter_203_io_enable = dut_io_coverage_102; // @[coverage.scala 106:31]
  assign SaturatingCounter_204_clock = clock;
  assign SaturatingCounter_204_reset = reset;
  assign SaturatingCounter_204_io_enable = ~dut_io_coverage_102; // @[coverage.scala 108:31]
  assign SaturatingCounter_205_clock = clock;
  assign SaturatingCounter_205_reset = reset;
  assign SaturatingCounter_205_io_enable = dut_io_coverage_103; // @[coverage.scala 106:31]
  assign SaturatingCounter_206_clock = clock;
  assign SaturatingCounter_206_reset = reset;
  assign SaturatingCounter_206_io_enable = ~dut_io_coverage_103; // @[coverage.scala 108:31]
  assign SaturatingCounter_207_clock = clock;
  assign SaturatingCounter_207_reset = reset;
  assign SaturatingCounter_207_io_enable = dut_io_coverage_104; // @[coverage.scala 106:31]
  assign SaturatingCounter_208_clock = clock;
  assign SaturatingCounter_208_reset = reset;
  assign SaturatingCounter_208_io_enable = ~dut_io_coverage_104; // @[coverage.scala 108:31]
  assign SaturatingCounter_209_clock = clock;
  assign SaturatingCounter_209_reset = reset;
  assign SaturatingCounter_209_io_enable = dut_io_coverage_105; // @[coverage.scala 106:31]
  assign SaturatingCounter_210_clock = clock;
  assign SaturatingCounter_210_reset = reset;
  assign SaturatingCounter_210_io_enable = ~dut_io_coverage_105; // @[coverage.scala 108:31]
  assign SaturatingCounter_211_clock = clock;
  assign SaturatingCounter_211_reset = reset;
  assign SaturatingCounter_211_io_enable = dut_io_coverage_106; // @[coverage.scala 106:31]
  assign SaturatingCounter_212_clock = clock;
  assign SaturatingCounter_212_reset = reset;
  assign SaturatingCounter_212_io_enable = ~dut_io_coverage_106; // @[coverage.scala 108:31]
  assign SaturatingCounter_213_clock = clock;
  assign SaturatingCounter_213_reset = reset;
  assign SaturatingCounter_213_io_enable = dut_io_coverage_107; // @[coverage.scala 106:31]
  assign SaturatingCounter_214_clock = clock;
  assign SaturatingCounter_214_reset = reset;
  assign SaturatingCounter_214_io_enable = ~dut_io_coverage_107; // @[coverage.scala 108:31]
  assign SaturatingCounter_215_clock = clock;
  assign SaturatingCounter_215_reset = reset;
  assign SaturatingCounter_215_io_enable = dut_io_coverage_108; // @[coverage.scala 106:31]
  assign SaturatingCounter_216_clock = clock;
  assign SaturatingCounter_216_reset = reset;
  assign SaturatingCounter_216_io_enable = ~dut_io_coverage_108; // @[coverage.scala 108:31]
  assign SaturatingCounter_217_clock = clock;
  assign SaturatingCounter_217_reset = reset;
  assign SaturatingCounter_217_io_enable = dut_io_coverage_109; // @[coverage.scala 106:31]
  assign SaturatingCounter_218_clock = clock;
  assign SaturatingCounter_218_reset = reset;
  assign SaturatingCounter_218_io_enable = ~dut_io_coverage_109; // @[coverage.scala 108:31]
  assign SaturatingCounter_219_clock = clock;
  assign SaturatingCounter_219_reset = reset;
  assign SaturatingCounter_219_io_enable = dut_io_coverage_110; // @[coverage.scala 106:31]
  assign SaturatingCounter_220_clock = clock;
  assign SaturatingCounter_220_reset = reset;
  assign SaturatingCounter_220_io_enable = ~dut_io_coverage_110; // @[coverage.scala 108:31]
  assign SaturatingCounter_221_clock = clock;
  assign SaturatingCounter_221_reset = reset;
  assign SaturatingCounter_221_io_enable = dut_io_coverage_111; // @[coverage.scala 106:31]
  assign SaturatingCounter_222_clock = clock;
  assign SaturatingCounter_222_reset = reset;
  assign SaturatingCounter_222_io_enable = ~dut_io_coverage_111; // @[coverage.scala 108:31]
  assign SaturatingCounter_223_clock = clock;
  assign SaturatingCounter_223_reset = reset;
  assign SaturatingCounter_223_io_enable = dut_io_coverage_112; // @[coverage.scala 106:31]
  assign SaturatingCounter_224_clock = clock;
  assign SaturatingCounter_224_reset = reset;
  assign SaturatingCounter_224_io_enable = ~dut_io_coverage_112; // @[coverage.scala 108:31]
  assign SaturatingCounter_225_clock = clock;
  assign SaturatingCounter_225_reset = reset;
  assign SaturatingCounter_225_io_enable = dut_io_coverage_113; // @[coverage.scala 106:31]
  assign SaturatingCounter_226_clock = clock;
  assign SaturatingCounter_226_reset = reset;
  assign SaturatingCounter_226_io_enable = ~dut_io_coverage_113; // @[coverage.scala 108:31]
  assign SaturatingCounter_227_clock = clock;
  assign SaturatingCounter_227_reset = reset;
  assign SaturatingCounter_227_io_enable = dut_io_coverage_114; // @[coverage.scala 106:31]
  assign SaturatingCounter_228_clock = clock;
  assign SaturatingCounter_228_reset = reset;
  assign SaturatingCounter_228_io_enable = ~dut_io_coverage_114; // @[coverage.scala 108:31]
  assign SaturatingCounter_229_clock = clock;
  assign SaturatingCounter_229_reset = reset;
  assign SaturatingCounter_229_io_enable = dut_io_coverage_115; // @[coverage.scala 106:31]
  assign SaturatingCounter_230_clock = clock;
  assign SaturatingCounter_230_reset = reset;
  assign SaturatingCounter_230_io_enable = ~dut_io_coverage_115; // @[coverage.scala 108:31]
  assign SaturatingCounter_231_clock = clock;
  assign SaturatingCounter_231_reset = reset;
  assign SaturatingCounter_231_io_enable = dut_io_coverage_116; // @[coverage.scala 106:31]
  assign SaturatingCounter_232_clock = clock;
  assign SaturatingCounter_232_reset = reset;
  assign SaturatingCounter_232_io_enable = ~dut_io_coverage_116; // @[coverage.scala 108:31]
  assign SaturatingCounter_233_clock = clock;
  assign SaturatingCounter_233_reset = reset;
  assign SaturatingCounter_233_io_enable = dut_io_coverage_117; // @[coverage.scala 106:31]
  assign SaturatingCounter_234_clock = clock;
  assign SaturatingCounter_234_reset = reset;
  assign SaturatingCounter_234_io_enable = ~dut_io_coverage_117; // @[coverage.scala 108:31]
  assign SaturatingCounter_235_clock = clock;
  assign SaturatingCounter_235_reset = reset;
  assign SaturatingCounter_235_io_enable = dut_io_coverage_118; // @[coverage.scala 106:31]
  assign SaturatingCounter_236_clock = clock;
  assign SaturatingCounter_236_reset = reset;
  assign SaturatingCounter_236_io_enable = ~dut_io_coverage_118; // @[coverage.scala 108:31]
  assign SaturatingCounter_237_clock = clock;
  assign SaturatingCounter_237_reset = reset;
  assign SaturatingCounter_237_io_enable = dut_io_coverage_119; // @[coverage.scala 106:31]
  assign SaturatingCounter_238_clock = clock;
  assign SaturatingCounter_238_reset = reset;
  assign SaturatingCounter_238_io_enable = ~dut_io_coverage_119; // @[coverage.scala 108:31]
  assign SaturatingCounter_239_clock = clock;
  assign SaturatingCounter_239_reset = reset;
  assign SaturatingCounter_239_io_enable = dut_io_coverage_120; // @[coverage.scala 106:31]
  assign SaturatingCounter_240_clock = clock;
  assign SaturatingCounter_240_reset = reset;
  assign SaturatingCounter_240_io_enable = ~dut_io_coverage_120; // @[coverage.scala 108:31]
  assign SaturatingCounter_241_clock = clock;
  assign SaturatingCounter_241_reset = reset;
  assign SaturatingCounter_241_io_enable = dut_io_coverage_121; // @[coverage.scala 106:31]
  assign SaturatingCounter_242_clock = clock;
  assign SaturatingCounter_242_reset = reset;
  assign SaturatingCounter_242_io_enable = ~dut_io_coverage_121; // @[coverage.scala 108:31]
  assign SaturatingCounter_243_clock = clock;
  assign SaturatingCounter_243_reset = reset;
  assign SaturatingCounter_243_io_enable = dut_io_coverage_122; // @[coverage.scala 106:31]
  assign SaturatingCounter_244_clock = clock;
  assign SaturatingCounter_244_reset = reset;
  assign SaturatingCounter_244_io_enable = ~dut_io_coverage_122; // @[coverage.scala 108:31]
  assign SaturatingCounter_245_clock = clock;
  assign SaturatingCounter_245_reset = reset;
  assign SaturatingCounter_245_io_enable = dut_io_coverage_123; // @[coverage.scala 106:31]
  assign SaturatingCounter_246_clock = clock;
  assign SaturatingCounter_246_reset = reset;
  assign SaturatingCounter_246_io_enable = ~dut_io_coverage_123; // @[coverage.scala 108:31]
  assign SaturatingCounter_247_clock = clock;
  assign SaturatingCounter_247_reset = reset;
  assign SaturatingCounter_247_io_enable = dut_io_coverage_124; // @[coverage.scala 106:31]
  assign SaturatingCounter_248_clock = clock;
  assign SaturatingCounter_248_reset = reset;
  assign SaturatingCounter_248_io_enable = ~dut_io_coverage_124; // @[coverage.scala 108:31]
  assign SaturatingCounter_249_clock = clock;
  assign SaturatingCounter_249_reset = reset;
  assign SaturatingCounter_249_io_enable = dut_io_coverage_125; // @[coverage.scala 106:31]
  assign SaturatingCounter_250_clock = clock;
  assign SaturatingCounter_250_reset = reset;
  assign SaturatingCounter_250_io_enable = ~dut_io_coverage_125; // @[coverage.scala 108:31]
  assign SaturatingCounter_251_clock = clock;
  assign SaturatingCounter_251_reset = reset;
  assign SaturatingCounter_251_io_enable = dut_io_coverage_126; // @[coverage.scala 106:31]
  assign SaturatingCounter_252_clock = clock;
  assign SaturatingCounter_252_reset = reset;
  assign SaturatingCounter_252_io_enable = ~dut_io_coverage_126; // @[coverage.scala 108:31]
  assign SaturatingCounter_253_clock = clock;
  assign SaturatingCounter_253_reset = reset;
  assign SaturatingCounter_253_io_enable = dut_io_coverage_127; // @[coverage.scala 106:31]
  assign SaturatingCounter_254_clock = clock;
  assign SaturatingCounter_254_reset = reset;
  assign SaturatingCounter_254_io_enable = ~dut_io_coverage_127; // @[coverage.scala 108:31]
  assign SaturatingCounter_255_clock = clock;
  assign SaturatingCounter_255_reset = reset;
  assign SaturatingCounter_255_io_enable = dut_io_coverage_128; // @[coverage.scala 106:31]
  assign SaturatingCounter_256_clock = clock;
  assign SaturatingCounter_256_reset = reset;
  assign SaturatingCounter_256_io_enable = ~dut_io_coverage_128; // @[coverage.scala 108:31]
  assign SaturatingCounter_257_clock = clock;
  assign SaturatingCounter_257_reset = reset;
  assign SaturatingCounter_257_io_enable = dut_io_coverage_129; // @[coverage.scala 106:31]
  assign SaturatingCounter_258_clock = clock;
  assign SaturatingCounter_258_reset = reset;
  assign SaturatingCounter_258_io_enable = ~dut_io_coverage_129; // @[coverage.scala 108:31]
  assign SaturatingCounter_259_clock = clock;
  assign SaturatingCounter_259_reset = reset;
  assign SaturatingCounter_259_io_enable = dut_io_coverage_130; // @[coverage.scala 106:31]
  assign SaturatingCounter_260_clock = clock;
  assign SaturatingCounter_260_reset = reset;
  assign SaturatingCounter_260_io_enable = ~dut_io_coverage_130; // @[coverage.scala 108:31]
  assign SaturatingCounter_261_clock = clock;
  assign SaturatingCounter_261_reset = reset;
  assign SaturatingCounter_261_io_enable = dut_io_coverage_131; // @[coverage.scala 106:31]
  assign SaturatingCounter_262_clock = clock;
  assign SaturatingCounter_262_reset = reset;
  assign SaturatingCounter_262_io_enable = ~dut_io_coverage_131; // @[coverage.scala 108:31]
  assign SaturatingCounter_263_clock = clock;
  assign SaturatingCounter_263_reset = reset;
  assign SaturatingCounter_263_io_enable = dut_io_coverage_132; // @[coverage.scala 106:31]
  assign SaturatingCounter_264_clock = clock;
  assign SaturatingCounter_264_reset = reset;
  assign SaturatingCounter_264_io_enable = ~dut_io_coverage_132; // @[coverage.scala 108:31]
  assign SaturatingCounter_265_clock = clock;
  assign SaturatingCounter_265_reset = reset;
  assign SaturatingCounter_265_io_enable = dut_io_coverage_133; // @[coverage.scala 106:31]
  assign SaturatingCounter_266_clock = clock;
  assign SaturatingCounter_266_reset = reset;
  assign SaturatingCounter_266_io_enable = ~dut_io_coverage_133; // @[coverage.scala 108:31]
  assign SaturatingCounter_267_clock = clock;
  assign SaturatingCounter_267_reset = reset;
  assign SaturatingCounter_267_io_enable = dut_io_coverage_134; // @[coverage.scala 106:31]
  assign SaturatingCounter_268_clock = clock;
  assign SaturatingCounter_268_reset = reset;
  assign SaturatingCounter_268_io_enable = ~dut_io_coverage_134; // @[coverage.scala 108:31]
  assign SaturatingCounter_269_clock = clock;
  assign SaturatingCounter_269_reset = reset;
  assign SaturatingCounter_269_io_enable = dut_io_coverage_135; // @[coverage.scala 106:31]
  assign SaturatingCounter_270_clock = clock;
  assign SaturatingCounter_270_reset = reset;
  assign SaturatingCounter_270_io_enable = ~dut_io_coverage_135; // @[coverage.scala 108:31]
  assign SaturatingCounter_271_clock = clock;
  assign SaturatingCounter_271_reset = reset;
  assign SaturatingCounter_271_io_enable = dut_io_coverage_136; // @[coverage.scala 106:31]
  assign SaturatingCounter_272_clock = clock;
  assign SaturatingCounter_272_reset = reset;
  assign SaturatingCounter_272_io_enable = ~dut_io_coverage_136; // @[coverage.scala 108:31]
  assign SaturatingCounter_273_clock = clock;
  assign SaturatingCounter_273_reset = reset;
  assign SaturatingCounter_273_io_enable = dut_io_coverage_137; // @[coverage.scala 106:31]
  assign SaturatingCounter_274_clock = clock;
  assign SaturatingCounter_274_reset = reset;
  assign SaturatingCounter_274_io_enable = ~dut_io_coverage_137; // @[coverage.scala 108:31]
  assign SaturatingCounter_275_clock = clock;
  assign SaturatingCounter_275_reset = reset;
  assign SaturatingCounter_275_io_enable = dut_io_coverage_138; // @[coverage.scala 106:31]
  assign SaturatingCounter_276_clock = clock;
  assign SaturatingCounter_276_reset = reset;
  assign SaturatingCounter_276_io_enable = ~dut_io_coverage_138; // @[coverage.scala 108:31]
  assign SaturatingCounter_277_clock = clock;
  assign SaturatingCounter_277_reset = reset;
  assign SaturatingCounter_277_io_enable = dut_io_coverage_139; // @[coverage.scala 106:31]
  assign SaturatingCounter_278_clock = clock;
  assign SaturatingCounter_278_reset = reset;
  assign SaturatingCounter_278_io_enable = ~dut_io_coverage_139; // @[coverage.scala 108:31]
  assign SaturatingCounter_279_clock = clock;
  assign SaturatingCounter_279_reset = reset;
  assign SaturatingCounter_279_io_enable = dut_io_coverage_140; // @[coverage.scala 106:31]
  assign SaturatingCounter_280_clock = clock;
  assign SaturatingCounter_280_reset = reset;
  assign SaturatingCounter_280_io_enable = ~dut_io_coverage_140; // @[coverage.scala 108:31]
  assign SaturatingCounter_281_clock = clock;
  assign SaturatingCounter_281_reset = reset;
  assign SaturatingCounter_281_io_enable = dut_io_coverage_141; // @[coverage.scala 106:31]
  assign SaturatingCounter_282_clock = clock;
  assign SaturatingCounter_282_reset = reset;
  assign SaturatingCounter_282_io_enable = ~dut_io_coverage_141; // @[coverage.scala 108:31]
  assign SaturatingCounter_283_clock = clock;
  assign SaturatingCounter_283_reset = reset;
  assign SaturatingCounter_283_io_enable = dut_io_coverage_142; // @[coverage.scala 106:31]
  assign SaturatingCounter_284_clock = clock;
  assign SaturatingCounter_284_reset = reset;
  assign SaturatingCounter_284_io_enable = ~dut_io_coverage_142; // @[coverage.scala 108:31]
  assign SaturatingCounter_285_clock = clock;
  assign SaturatingCounter_285_reset = reset;
  assign SaturatingCounter_285_io_enable = dut_io_coverage_143; // @[coverage.scala 106:31]
  assign SaturatingCounter_286_clock = clock;
  assign SaturatingCounter_286_reset = reset;
  assign SaturatingCounter_286_io_enable = ~dut_io_coverage_143; // @[coverage.scala 108:31]
  assign SaturatingCounter_287_clock = clock;
  assign SaturatingCounter_287_reset = reset;
  assign SaturatingCounter_287_io_enable = dut_io_coverage_144; // @[coverage.scala 106:31]
  assign SaturatingCounter_288_clock = clock;
  assign SaturatingCounter_288_reset = reset;
  assign SaturatingCounter_288_io_enable = ~dut_io_coverage_144; // @[coverage.scala 108:31]
  assign SaturatingCounter_289_clock = clock;
  assign SaturatingCounter_289_reset = reset;
  assign SaturatingCounter_289_io_enable = dut_io_coverage_145; // @[coverage.scala 106:31]
  assign SaturatingCounter_290_clock = clock;
  assign SaturatingCounter_290_reset = reset;
  assign SaturatingCounter_290_io_enable = ~dut_io_coverage_145; // @[coverage.scala 108:31]
  assign SaturatingCounter_291_clock = clock;
  assign SaturatingCounter_291_reset = reset;
  assign SaturatingCounter_291_io_enable = dut_io_coverage_146; // @[coverage.scala 106:31]
  assign SaturatingCounter_292_clock = clock;
  assign SaturatingCounter_292_reset = reset;
  assign SaturatingCounter_292_io_enable = ~dut_io_coverage_146; // @[coverage.scala 108:31]
  assign SaturatingCounter_293_clock = clock;
  assign SaturatingCounter_293_reset = reset;
  assign SaturatingCounter_293_io_enable = dut_io_coverage_147; // @[coverage.scala 106:31]
  assign SaturatingCounter_294_clock = clock;
  assign SaturatingCounter_294_reset = reset;
  assign SaturatingCounter_294_io_enable = ~dut_io_coverage_147; // @[coverage.scala 108:31]
  assign SaturatingCounter_295_clock = clock;
  assign SaturatingCounter_295_reset = reset;
  assign SaturatingCounter_295_io_enable = dut_io_coverage_148; // @[coverage.scala 106:31]
  assign SaturatingCounter_296_clock = clock;
  assign SaturatingCounter_296_reset = reset;
  assign SaturatingCounter_296_io_enable = ~dut_io_coverage_148; // @[coverage.scala 108:31]
  assign SaturatingCounter_297_clock = clock;
  assign SaturatingCounter_297_reset = reset;
  assign SaturatingCounter_297_io_enable = dut_io_coverage_149; // @[coverage.scala 106:31]
  assign SaturatingCounter_298_clock = clock;
  assign SaturatingCounter_298_reset = reset;
  assign SaturatingCounter_298_io_enable = ~dut_io_coverage_149; // @[coverage.scala 108:31]
  assign SaturatingCounter_299_clock = clock;
  assign SaturatingCounter_299_reset = reset;
  assign SaturatingCounter_299_io_enable = dut_io_coverage_150; // @[coverage.scala 106:31]
  assign SaturatingCounter_300_clock = clock;
  assign SaturatingCounter_300_reset = reset;
  assign SaturatingCounter_300_io_enable = ~dut_io_coverage_150; // @[coverage.scala 108:31]
  assign SaturatingCounter_301_clock = clock;
  assign SaturatingCounter_301_reset = reset;
  assign SaturatingCounter_301_io_enable = dut_io_coverage_151; // @[coverage.scala 106:31]
  assign SaturatingCounter_302_clock = clock;
  assign SaturatingCounter_302_reset = reset;
  assign SaturatingCounter_302_io_enable = ~dut_io_coverage_151; // @[coverage.scala 108:31]
  assign SaturatingCounter_303_clock = clock;
  assign SaturatingCounter_303_reset = reset;
  assign SaturatingCounter_303_io_enable = dut_io_coverage_152; // @[coverage.scala 106:31]
  assign SaturatingCounter_304_clock = clock;
  assign SaturatingCounter_304_reset = reset;
  assign SaturatingCounter_304_io_enable = ~dut_io_coverage_152; // @[coverage.scala 108:31]
  assign SaturatingCounter_305_clock = clock;
  assign SaturatingCounter_305_reset = reset;
  assign SaturatingCounter_305_io_enable = dut_io_coverage_153; // @[coverage.scala 106:31]
  assign SaturatingCounter_306_clock = clock;
  assign SaturatingCounter_306_reset = reset;
  assign SaturatingCounter_306_io_enable = ~dut_io_coverage_153; // @[coverage.scala 108:31]
  assign SaturatingCounter_307_clock = clock;
  assign SaturatingCounter_307_reset = reset;
  assign SaturatingCounter_307_io_enable = dut_io_coverage_154; // @[coverage.scala 106:31]
  assign SaturatingCounter_308_clock = clock;
  assign SaturatingCounter_308_reset = reset;
  assign SaturatingCounter_308_io_enable = ~dut_io_coverage_154; // @[coverage.scala 108:31]
  assign SaturatingCounter_309_clock = clock;
  assign SaturatingCounter_309_reset = reset;
  assign SaturatingCounter_309_io_enable = dut_io_coverage_155; // @[coverage.scala 106:31]
  assign SaturatingCounter_310_clock = clock;
  assign SaturatingCounter_310_reset = reset;
  assign SaturatingCounter_310_io_enable = ~dut_io_coverage_155; // @[coverage.scala 108:31]
  assign SaturatingCounter_311_clock = clock;
  assign SaturatingCounter_311_reset = reset;
  assign SaturatingCounter_311_io_enable = dut_io_coverage_156; // @[coverage.scala 106:31]
  assign SaturatingCounter_312_clock = clock;
  assign SaturatingCounter_312_reset = reset;
  assign SaturatingCounter_312_io_enable = ~dut_io_coverage_156; // @[coverage.scala 108:31]
  assign SaturatingCounter_313_clock = clock;
  assign SaturatingCounter_313_reset = reset;
  assign SaturatingCounter_313_io_enable = dut_io_coverage_157; // @[coverage.scala 106:31]
  assign SaturatingCounter_314_clock = clock;
  assign SaturatingCounter_314_reset = reset;
  assign SaturatingCounter_314_io_enable = ~dut_io_coverage_157; // @[coverage.scala 108:31]
  assign SaturatingCounter_315_clock = clock;
  assign SaturatingCounter_315_reset = reset;
  assign SaturatingCounter_315_io_enable = dut_io_coverage_158; // @[coverage.scala 106:31]
  assign SaturatingCounter_316_clock = clock;
  assign SaturatingCounter_316_reset = reset;
  assign SaturatingCounter_316_io_enable = ~dut_io_coverage_158; // @[coverage.scala 108:31]
  assign SaturatingCounter_317_clock = clock;
  assign SaturatingCounter_317_reset = reset;
  assign SaturatingCounter_317_io_enable = dut_io_coverage_159; // @[coverage.scala 106:31]
  assign SaturatingCounter_318_clock = clock;
  assign SaturatingCounter_318_reset = reset;
  assign SaturatingCounter_318_io_enable = ~dut_io_coverage_159; // @[coverage.scala 108:31]
  assign SaturatingCounter_319_clock = clock;
  assign SaturatingCounter_319_reset = reset;
  assign SaturatingCounter_319_io_enable = dut_io_coverage_160; // @[coverage.scala 106:31]
  assign SaturatingCounter_320_clock = clock;
  assign SaturatingCounter_320_reset = reset;
  assign SaturatingCounter_320_io_enable = ~dut_io_coverage_160; // @[coverage.scala 108:31]
  assign SaturatingCounter_321_clock = clock;
  assign SaturatingCounter_321_reset = reset;
  assign SaturatingCounter_321_io_enable = dut_io_coverage_161; // @[coverage.scala 106:31]
  assign SaturatingCounter_322_clock = clock;
  assign SaturatingCounter_322_reset = reset;
  assign SaturatingCounter_322_io_enable = ~dut_io_coverage_161; // @[coverage.scala 108:31]
  assign SaturatingCounter_323_clock = clock;
  assign SaturatingCounter_323_reset = reset;
  assign SaturatingCounter_323_io_enable = dut_io_coverage_162; // @[coverage.scala 106:31]
  assign SaturatingCounter_324_clock = clock;
  assign SaturatingCounter_324_reset = reset;
  assign SaturatingCounter_324_io_enable = ~dut_io_coverage_162; // @[coverage.scala 108:31]
  assign SaturatingCounter_325_clock = clock;
  assign SaturatingCounter_325_reset = reset;
  assign SaturatingCounter_325_io_enable = dut_io_coverage_163; // @[coverage.scala 106:31]
  assign SaturatingCounter_326_clock = clock;
  assign SaturatingCounter_326_reset = reset;
  assign SaturatingCounter_326_io_enable = ~dut_io_coverage_163; // @[coverage.scala 108:31]
  assign SaturatingCounter_327_clock = clock;
  assign SaturatingCounter_327_reset = reset;
  assign SaturatingCounter_327_io_enable = dut_io_coverage_164; // @[coverage.scala 106:31]
  assign SaturatingCounter_328_clock = clock;
  assign SaturatingCounter_328_reset = reset;
  assign SaturatingCounter_328_io_enable = ~dut_io_coverage_164; // @[coverage.scala 108:31]
  assign SaturatingCounter_329_clock = clock;
  assign SaturatingCounter_329_reset = reset;
  assign SaturatingCounter_329_io_enable = dut_io_coverage_165; // @[coverage.scala 106:31]
  assign SaturatingCounter_330_clock = clock;
  assign SaturatingCounter_330_reset = reset;
  assign SaturatingCounter_330_io_enable = ~dut_io_coverage_165; // @[coverage.scala 108:31]
  assign SaturatingCounter_331_clock = clock;
  assign SaturatingCounter_331_reset = reset;
  assign SaturatingCounter_331_io_enable = dut_io_coverage_166; // @[coverage.scala 106:31]
  assign SaturatingCounter_332_clock = clock;
  assign SaturatingCounter_332_reset = reset;
  assign SaturatingCounter_332_io_enable = ~dut_io_coverage_166; // @[coverage.scala 108:31]
  assign SaturatingCounter_333_clock = clock;
  assign SaturatingCounter_333_reset = reset;
  assign SaturatingCounter_333_io_enable = dut_io_coverage_167; // @[coverage.scala 106:31]
  assign SaturatingCounter_334_clock = clock;
  assign SaturatingCounter_334_reset = reset;
  assign SaturatingCounter_334_io_enable = ~dut_io_coverage_167; // @[coverage.scala 108:31]
  assign SaturatingCounter_335_clock = clock;
  assign SaturatingCounter_335_reset = reset;
  assign SaturatingCounter_335_io_enable = dut_io_coverage_168; // @[coverage.scala 106:31]
  assign SaturatingCounter_336_clock = clock;
  assign SaturatingCounter_336_reset = reset;
  assign SaturatingCounter_336_io_enable = ~dut_io_coverage_168; // @[coverage.scala 108:31]
  assign SaturatingCounter_337_clock = clock;
  assign SaturatingCounter_337_reset = reset;
  assign SaturatingCounter_337_io_enable = dut_io_coverage_169; // @[coverage.scala 106:31]
  assign SaturatingCounter_338_clock = clock;
  assign SaturatingCounter_338_reset = reset;
  assign SaturatingCounter_338_io_enable = ~dut_io_coverage_169; // @[coverage.scala 108:31]
  assign SaturatingCounter_339_clock = clock;
  assign SaturatingCounter_339_reset = reset;
  assign SaturatingCounter_339_io_enable = dut_io_coverage_170; // @[coverage.scala 106:31]
  assign SaturatingCounter_340_clock = clock;
  assign SaturatingCounter_340_reset = reset;
  assign SaturatingCounter_340_io_enable = ~dut_io_coverage_170; // @[coverage.scala 108:31]
  assign SaturatingCounter_341_clock = clock;
  assign SaturatingCounter_341_reset = reset;
  assign SaturatingCounter_341_io_enable = dut_io_coverage_171; // @[coverage.scala 106:31]
  assign SaturatingCounter_342_clock = clock;
  assign SaturatingCounter_342_reset = reset;
  assign SaturatingCounter_342_io_enable = ~dut_io_coverage_171; // @[coverage.scala 108:31]
  assign SaturatingCounter_343_clock = clock;
  assign SaturatingCounter_343_reset = reset;
  assign SaturatingCounter_343_io_enable = dut_io_coverage_172; // @[coverage.scala 106:31]
  assign SaturatingCounter_344_clock = clock;
  assign SaturatingCounter_344_reset = reset;
  assign SaturatingCounter_344_io_enable = ~dut_io_coverage_172; // @[coverage.scala 108:31]
  assign SaturatingCounter_345_clock = clock;
  assign SaturatingCounter_345_reset = reset;
  assign SaturatingCounter_345_io_enable = dut_io_coverage_173; // @[coverage.scala 106:31]
  assign SaturatingCounter_346_clock = clock;
  assign SaturatingCounter_346_reset = reset;
  assign SaturatingCounter_346_io_enable = ~dut_io_coverage_173; // @[coverage.scala 108:31]
  assign SaturatingCounter_347_clock = clock;
  assign SaturatingCounter_347_reset = reset;
  assign SaturatingCounter_347_io_enable = dut_io_coverage_174; // @[coverage.scala 106:31]
  assign SaturatingCounter_348_clock = clock;
  assign SaturatingCounter_348_reset = reset;
  assign SaturatingCounter_348_io_enable = ~dut_io_coverage_174; // @[coverage.scala 108:31]
  assign SaturatingCounter_349_clock = clock;
  assign SaturatingCounter_349_reset = reset;
  assign SaturatingCounter_349_io_enable = dut_io_coverage_175; // @[coverage.scala 106:31]
  assign SaturatingCounter_350_clock = clock;
  assign SaturatingCounter_350_reset = reset;
  assign SaturatingCounter_350_io_enable = ~dut_io_coverage_175; // @[coverage.scala 108:31]
  assign SaturatingCounter_351_clock = clock;
  assign SaturatingCounter_351_reset = reset;
  assign SaturatingCounter_351_io_enable = dut_io_coverage_176; // @[coverage.scala 106:31]
  assign SaturatingCounter_352_clock = clock;
  assign SaturatingCounter_352_reset = reset;
  assign SaturatingCounter_352_io_enable = ~dut_io_coverage_176; // @[coverage.scala 108:31]
  assign SaturatingCounter_353_clock = clock;
  assign SaturatingCounter_353_reset = reset;
  assign SaturatingCounter_353_io_enable = dut_io_coverage_177; // @[coverage.scala 106:31]
  assign SaturatingCounter_354_clock = clock;
  assign SaturatingCounter_354_reset = reset;
  assign SaturatingCounter_354_io_enable = ~dut_io_coverage_177; // @[coverage.scala 108:31]
  assign SaturatingCounter_355_clock = clock;
  assign SaturatingCounter_355_reset = reset;
  assign SaturatingCounter_355_io_enable = dut_io_coverage_178; // @[coverage.scala 106:31]
  assign SaturatingCounter_356_clock = clock;
  assign SaturatingCounter_356_reset = reset;
  assign SaturatingCounter_356_io_enable = ~dut_io_coverage_178; // @[coverage.scala 108:31]
  assign SaturatingCounter_357_clock = clock;
  assign SaturatingCounter_357_reset = reset;
  assign SaturatingCounter_357_io_enable = dut_io_coverage_179; // @[coverage.scala 106:31]
  assign SaturatingCounter_358_clock = clock;
  assign SaturatingCounter_358_reset = reset;
  assign SaturatingCounter_358_io_enable = ~dut_io_coverage_179; // @[coverage.scala 108:31]
  assign SaturatingCounter_359_clock = clock;
  assign SaturatingCounter_359_reset = reset;
  assign SaturatingCounter_359_io_enable = dut_io_coverage_180; // @[coverage.scala 106:31]
  assign SaturatingCounter_360_clock = clock;
  assign SaturatingCounter_360_reset = reset;
  assign SaturatingCounter_360_io_enable = ~dut_io_coverage_180; // @[coverage.scala 108:31]
  assign SaturatingCounter_361_clock = clock;
  assign SaturatingCounter_361_reset = reset;
  assign SaturatingCounter_361_io_enable = dut_io_coverage_181; // @[coverage.scala 106:31]
  assign SaturatingCounter_362_clock = clock;
  assign SaturatingCounter_362_reset = reset;
  assign SaturatingCounter_362_io_enable = ~dut_io_coverage_181; // @[coverage.scala 108:31]
  assign SaturatingCounter_363_clock = clock;
  assign SaturatingCounter_363_reset = reset;
  assign SaturatingCounter_363_io_enable = dut_io_coverage_182; // @[coverage.scala 106:31]
  assign SaturatingCounter_364_clock = clock;
  assign SaturatingCounter_364_reset = reset;
  assign SaturatingCounter_364_io_enable = ~dut_io_coverage_182; // @[coverage.scala 108:31]
  assign SaturatingCounter_365_clock = clock;
  assign SaturatingCounter_365_reset = reset;
  assign SaturatingCounter_365_io_enable = dut_io_coverage_183; // @[coverage.scala 106:31]
  assign SaturatingCounter_366_clock = clock;
  assign SaturatingCounter_366_reset = reset;
  assign SaturatingCounter_366_io_enable = ~dut_io_coverage_183; // @[coverage.scala 108:31]
  assign SaturatingCounter_367_clock = clock;
  assign SaturatingCounter_367_reset = reset;
  assign SaturatingCounter_367_io_enable = dut_io_coverage_184; // @[coverage.scala 106:31]
  assign SaturatingCounter_368_clock = clock;
  assign SaturatingCounter_368_reset = reset;
  assign SaturatingCounter_368_io_enable = ~dut_io_coverage_184; // @[coverage.scala 108:31]
  assign SaturatingCounter_369_clock = clock;
  assign SaturatingCounter_369_reset = reset;
  assign SaturatingCounter_369_io_enable = dut_io_coverage_185; // @[coverage.scala 106:31]
  assign SaturatingCounter_370_clock = clock;
  assign SaturatingCounter_370_reset = reset;
  assign SaturatingCounter_370_io_enable = ~dut_io_coverage_185; // @[coverage.scala 108:31]
  assign SaturatingCounter_371_clock = clock;
  assign SaturatingCounter_371_reset = reset;
  assign SaturatingCounter_371_io_enable = dut_io_coverage_186; // @[coverage.scala 106:31]
  assign SaturatingCounter_372_clock = clock;
  assign SaturatingCounter_372_reset = reset;
  assign SaturatingCounter_372_io_enable = ~dut_io_coverage_186; // @[coverage.scala 108:31]
endmodule
