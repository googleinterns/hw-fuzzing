module Sodor3Stage(
  input          metaReset,
  input          clock,
  input          reset,
  input          io_imem_req_ready,
  output         io_imem_req_valid,
  output [31:0]  io_imem_req_bits_addr,
  output [31:0]  io_imem_req_bits_data,
  output         io_imem_req_bits_fcn,
  output [2:0]   io_imem_req_bits_typ,
  input          io_imem_resp_valid,
  input  [31:0]  io_imem_resp_bits_data,
  input          io_reset,
  output         assert_out,
  output [615:0] auto_cover_out
);
  wire  core_metaReset; // @[top.scala 26:26]
  wire  core_clock; // @[top.scala 26:26]
  wire  core_reset; // @[top.scala 26:26]
  wire [31:0] core_io_imem_req_bits_addr; // @[top.scala 26:26]
  wire [31:0] core_io_imem_resp_bits_data; // @[top.scala 26:26]
  wire [31:0] core_io_dmem_req_bits_addr; // @[top.scala 26:26]
  wire [31:0] core_io_dmem_req_bits_data; // @[top.scala 26:26]
  wire  core_io_dmem_req_bits_fcn; // @[top.scala 26:26]
  wire [2:0] core_io_dmem_req_bits_typ; // @[top.scala 26:26]
  wire [31:0] core_io_dmem_resp_bits_data; // @[top.scala 26:26]
  wire  core__GEN_411; // @[top.scala 26:26]
  wire  core__GEN_405; // @[top.scala 26:26]
  wire  core__GEN_92; // @[top.scala 26:26]
  wire  core__GEN_52; // @[top.scala 26:26]
  wire  core__GEN_305; // @[top.scala 26:26]
  wire  core__GEN_200; // @[top.scala 26:26]
  wire  core__GEN_149; // @[top.scala 26:26]
  wire  core__GEN_426; // @[top.scala 26:26]
  wire  core__GEN_291; // @[top.scala 26:26]
  wire  core__GEN_1_0; // @[top.scala 26:26]
  wire  core__GEN_25; // @[top.scala 26:26]
  wire  core__GEN_248; // @[top.scala 26:26]
  wire  core__GEN_107; // @[top.scala 26:26]
  wire  core__GEN_134; // @[top.scala 26:26]
  wire  core__GEN_206; // @[top.scala 26:26]
  wire  core__GEN_40; // @[top.scala 26:26]
  wire  core__GEN_306; // @[top.scala 26:26]
  wire  core__GEN_233; // @[top.scala 26:26]
  wire  core__GEN_128; // @[top.scala 26:26]
  wire  core__GEN_384; // @[top.scala 26:26]
  wire  core__GEN_191; // @[top.scala 26:26]
  wire  core__GEN_16; // @[top.scala 26:26]
  wire  core__GEN_227; // @[top.scala 26:26]
  wire  core__GEN_19; // @[top.scala 26:26]
  wire  core__GEN_327; // @[top.scala 26:26]
  wire  core__GEN_113; // @[top.scala 26:26]
  wire  core__GEN_46; // @[top.scala 26:26]
  wire  core__GEN_299; // @[top.scala 26:26]
  wire  core__GEN_390; // @[top.scala 26:26]
  wire  core__GEN_73; // @[top.scala 26:26]
  wire  core__GEN_212; // @[top.scala 26:26]
  wire  core__GEN_10; // @[top.scala 26:26]
  wire  core__GEN_285; // @[top.scala 26:26]
  wire  core__GEN_318; // @[top.scala 26:26]
  wire  core__GEN_312; // @[top.scala 26:26]
  wire  core__GEN_31; // @[top.scala 26:26]
  wire  core__GEN_311; // @[top.scala 26:26]
  wire  core__GEN_67; // @[top.scala 26:26]
  wire  core__GEN_320; // @[top.scala 26:26]
  wire  core__GEN_399; // @[top.scala 26:26]
  wire  core__GEN_215; // @[top.scala 26:26]
  wire  core__GEN_221; // @[top.scala 26:26]
  wire  core__GEN_101; // @[top.scala 26:26]
  wire  core__GEN_110; // @[top.scala 26:26]
  wire  core__GEN_387; // @[top.scala 26:26]
  wire  core__GEN_283; // @[top.scala 26:26]
  wire  core__GEN_314; // @[top.scala 26:26]
  wire  core__GEN_178; // @[top.scala 26:26]
  wire  core__GEN_209; // @[top.scala 26:26]
  wire  core__GEN_300; // @[top.scala 26:26]
  wire  core__GEN_279; // @[top.scala 26:26]
  wire  core__GEN_269; // @[top.scala 26:26]
  wire  core__GEN_28; // @[top.scala 26:26]
  wire  core__GEN_277; // @[top.scala 26:26]
  wire  core__GEN_378; // @[top.scala 26:26]
  wire  core__GEN_368; // @[top.scala 26:26]
  wire  core__GEN_55; // @[top.scala 26:26]
  wire  core__GEN_377; // @[top.scala 26:26]
  wire  core__GEN_194; // @[top.scala 26:26]
  wire  core__GEN_22; // @[top.scala 26:26]
  wire  core__GEN_12; // @[top.scala 26:26]
  wire  core__GEN_294; // @[top.scala 26:26]
  wire  core__GEN_13; // @[top.scala 26:26]
  wire  core__GEN_49; // @[top.scala 26:26]
  wire  core__GEN_116; // @[top.scala 26:26]
  wire  core__GEN_393; // @[top.scala 26:26]
  wire  core__GEN_362; // @[top.scala 26:26]
  wire  core__GEN_7; // @[top.scala 26:26]
  wire  core__GEN_461; // @[top.scala 26:26]
  wire  core__GEN_34; // @[top.scala 26:26]
  wire  core__GEN_122; // @[top.scala 26:26]
  wire  core__GEN_308; // @[top.scala 26:26]
  wire  core__GEN_263; // @[top.scala 26:26]
  wire  core__GEN_95; // @[top.scala 26:26]
  wire  core__GEN_230; // @[top.scala 26:26]
  wire  core__GEN_293; // @[top.scala 26:26]
  wire  core__GEN_184; // @[top.scala 26:26]
  wire  core__GEN_1_1; // @[top.scala 26:26]
  wire  core__GEN_10_0; // @[top.scala 26:26]
  wire  core__GEN_197; // @[top.scala 26:26]
  wire  core__GEN_187; // @[top.scala 26:26]
  wire  core__GEN_449; // @[top.scala 26:26]
  wire  core__GEN_288; // @[top.scala 26:26]
  wire  core__GEN_104; // @[top.scala 26:26]
  wire  core__GEN_265; // @[top.scala 26:26]
  wire  core__GEN_296; // @[top.scala 26:26]
  wire  core__GEN_160; // @[top.scala 26:26]
  wire  core__GEN_172; // @[top.scala 26:26]
  wire  core__GEN_203; // @[top.scala 26:26]
  wire  core__GEN_245; // @[top.scala 26:26]
  wire  core__GEN_0; // @[top.scala 26:26]
  wire  core__GEN_272; // @[top.scala 26:26]
  wire  core__GEN_271; // @[top.scala 26:26]
  wire  core__GEN_37; // @[top.scala 26:26]
  wire  core__GEN_166; // @[top.scala 26:26]
  wire  core__GEN_280; // @[top.scala 26:26]
  wire  core__GEN_286; // @[top.scala 26:26]
  wire  core__GEN_381; // @[top.scala 26:26]
  wire  core__GEN_371; // @[top.scala 26:26]
  wire  core__GEN_266; // @[top.scala 26:26]
  wire  core__GEN_16_0; // @[top.scala 26:26]
  wire  core__GEN_22_0; // @[top.scala 26:26]
  wire  core__GEN_302; // @[top.scala 26:26]
  wire  core__GEN_344; // @[top.scala 26:26]
  wire  core__GEN_282; // @[top.scala 26:26]
  wire  core__GEN_443; // @[top.scala 26:26]
  wire  core__GEN_16_1; // @[top.scala 26:26]
  wire  core__GEN_251; // @[top.scala 26:26]
  wire  core__GEN_10_1; // @[top.scala 26:26]
  wire  core__GEN_259; // @[top.scala 26:26]
  wire  core__GEN_98; // @[top.scala 26:26]
  wire  core__GEN_6; // @[top.scala 26:26]
  wire  core__GEN_350; // @[top.scala 26:26]
  wire  core__GEN_365; // @[top.scala 26:26]
  wire  core__GEN_15; // @[top.scala 26:26]
  wire  core__GEN_152; // @[top.scala 26:26]
  wire  core__GEN_446; // @[top.scala 26:26]
  wire  core__GEN_332; // @[top.scala 26:26]
  wire  core__GEN_326; // @[top.scala 26:26]
  wire  core__GEN_19_0; // @[top.scala 26:26]
  wire  core__GEN_148; // @[top.scala 26:26]
  wire  core__GEN_359; // @[top.scala 26:26]
  wire  core__GEN_15_0; // @[top.scala 26:26]
  wire  core__GEN_87; // @[top.scala 26:26]
  wire  core__GEN_458; // @[top.scala 26:26]
  wire  core__GEN_452; // @[top.scala 26:26]
  wire  core__GEN_13_0; // @[top.scala 26:26]
  wire  core__GEN_3; // @[top.scala 26:26]
  wire  core__GEN_347; // @[top.scala 26:26]
  wire  core__GEN_274; // @[top.scala 26:26]
  wire  core__GEN_425; // @[top.scala 26:26]
  wire  core__GEN_239; // @[top.scala 26:26]
  wire  core__GEN_232; // @[top.scala 26:26]
  wire  core__GEN_190; // @[top.scala 26:26]
  wire  core__GEN_154; // @[top.scala 26:26]
  wire  core__GEN_289; // @[top.scala 26:26]
  wire  core__GEN_431; // @[top.scala 26:26]
  wire  core__GEN_181; // @[top.scala 26:26]
  wire  core__GEN_253; // @[top.scala 26:26]
  wire  core__GEN_254; // @[top.scala 26:26]
  wire  core__GEN_353; // @[top.scala 26:26]
  wire  core__GEN_72; // @[top.scala 26:26]
  wire  core__GEN_175; // @[top.scala 26:26]
  wire  core__GEN_169; // @[top.scala 26:26]
  wire  core__GEN_260; // @[top.scala 26:26]
  wire  core__GEN_4_0; // @[top.scala 26:26]
  wire  core__GEN_275; // @[top.scala 26:26]
  wire  core__GEN_247; // @[top.scala 26:26]
  wire  core__GEN_268; // @[top.scala 26:26]
  wire  core__GEN_9; // @[top.scala 26:26]
  wire  core__GEN_338; // @[top.scala 26:26]
  wire  core__GEN_374; // @[top.scala 26:26]
  wire  core__GEN_242; // @[top.scala 26:26]
  wire  core__GEN_214; // @[top.scala 26:26]
  wire  core__GEN_250; // @[top.scala 26:26]
  wire  core__GEN_455; // @[top.scala 26:26]
  wire  core__GEN_241; // @[top.scala 26:26]
  wire  core__GEN_142; // @[top.scala 26:26]
  wire  core__GEN_136; // @[top.scala 26:26]
  wire  core__GEN_413; // @[top.scala 26:26]
  wire  core__GEN_235; // @[top.scala 26:26]
  wire  core__GEN_236; // @[top.scala 26:26]
  wire  core__GEN_262; // @[top.scala 26:26]
  wire  core__GEN_335; // @[top.scala 26:26]
  wire  core__GEN_54; // @[top.scala 26:26]
  wire  core__GEN_313; // @[top.scala 26:26]
  wire  core__GEN_18; // @[top.scala 26:26]
  wire  core__GEN_69; // @[top.scala 26:26]
  wire  core__GEN_157; // @[top.scala 26:26]
  wire  core__GEN_434; // @[top.scala 26:26]
  wire  core__GEN_248_0; // @[top.scala 26:26]
  wire  core__GEN_257; // @[top.scala 26:26]
  wire  core__GEN_320_0; // @[top.scala 26:26]
  wire  core__GEN_75; // @[top.scala 26:26]
  wire  core__GEN_356; // @[top.scala 26:26]
  wire  core__GEN_12_0; // @[top.scala 26:26]
  wire  core__GEN_90; // @[top.scala 26:26]
  wire  core__GEN_163; // @[top.scala 26:26]
  wire  core__GEN_419; // @[top.scala 26:26]
  wire  core__GEN_314_0; // @[top.scala 26:26]
  wire  core__GEN_7_0; // @[top.scala 26:26]
  wire  core__GEN_130; // @[top.scala 26:26]
  wire  core__GEN_341; // @[top.scala 26:26]
  wire  core__GEN_440; // @[top.scala 26:26]
  wire  core__GEN_229; // @[top.scala 26:26]
  wire  core__GEN_299_0; // @[top.scala 26:26]
  wire  core__GEN_121; // @[top.scala 26:26]
  wire  core__GEN_256; // @[top.scala 26:26]
  wire  core__GEN_398; // @[top.scala 26:26]
  wire  core__GEN_81; // @[top.scala 26:26]
  wire  core__GEN_407; // @[top.scala 26:26]
  wire  core__GEN_149_0; // @[top.scala 26:26]
  wire  core__GEN_416; // @[top.scala 26:26]
  wire  core__GEN_281; // @[top.scala 26:26]
  wire  core__GEN_15_1; // @[top.scala 26:26]
  wire  core__GEN_380; // @[top.scala 26:26]
  wire  core__GEN_57; // @[top.scala 26:26]
  wire  core__GEN_145; // @[top.scala 26:26]
  wire  core__GEN_296_0; // @[top.scala 26:26]
  wire  core__GEN_223; // @[top.scala 26:26]
  wire  core__GEN_118; // @[top.scala 26:26]
  wire  core__GEN_322; // @[top.scala 26:26]
  wire  core__GEN_422; // @[top.scala 26:26]
  wire  core__GEN_244; // @[top.scala 26:26]
  wire  core__GEN_124; // @[top.scala 26:26]
  wire  core__GEN_103; // @[top.scala 26:26]
  wire  core__GEN_238; // @[top.scala 26:26]
  wire  core__GEN_329; // @[top.scala 26:26]
  wire  core__GEN_63; // @[top.scala 26:26]
  wire  core__GEN_151; // @[top.scala 26:26]
  wire  core__GEN_202; // @[top.scala 26:26]
  wire  core__GEN_6_0; // @[top.scala 26:26]
  wire  core__GEN_196; // @[top.scala 26:26]
  wire  core__GEN_437; // @[top.scala 26:26]
  wire  core__GEN_302_0; // @[top.scala 26:26]
  wire  core__GEN_295; // @[top.scala 26:26]
  wire  core__GEN_301; // @[top.scala 26:26]
  wire  core__GEN_310; // @[top.scala 26:26]
  wire  core__GEN_401; // @[top.scala 26:26]
  wire  core__GEN_395; // @[top.scala 26:26]
  wire  core__GEN_78; // @[top.scala 26:26]
  wire  core__GEN_84; // @[top.scala 26:26]
  wire  core__GEN_217; // @[top.scala 26:26]
  wire  core__GEN_428; // @[top.scala 26:26]
  wire  core__GEN_308_0; // @[top.scala 26:26]
  wire  core__GEN_323; // @[top.scala 26:26]
  wire  core__GEN_36; // @[top.scala 26:26]
  wire  core__GEN_42; // @[top.scala 26:26]
  wire  core__GEN_317; // @[top.scala 26:26]
  wire  core__GEN_316; // @[top.scala 26:26]
  wire  core__GEN_139; // @[top.scala 26:26]
  wire  core__GEN_404; // @[top.scala 26:26]
  wire  core__GEN_290; // @[top.scala 26:26]
  wire  core__GEN_18_0; // @[top.scala 26:26]
  wire  core__GEN_226; // @[top.scala 26:26]
  wire  core__GEN_106; // @[top.scala 26:26]
  wire  core__GEN_51; // @[top.scala 26:26]
  wire  core__GEN_45; // @[top.scala 26:26]
  wire  core__GEN_9_0; // @[top.scala 26:26]
  wire  core__GEN_367; // @[top.scala 26:26]
  wire  core__GEN_319; // @[top.scala 26:26]
  wire  core__GEN_284; // @[top.scala 26:26]
  wire  core__GEN_274_0; // @[top.scala 26:26]
  wire  core__GEN_39; // @[top.scala 26:26]
  wire  core__GEN_383; // @[top.scala 26:26]
  wire  core__GEN_373; // @[top.scala 26:26]
  wire  core__GEN_66; // @[top.scala 26:26]
  wire  core__GEN_18_1; // @[top.scala 26:26]
  wire  core__GEN_410; // @[top.scala 26:26]
  wire  core__GEN_24; // @[top.scala 26:26]
  wire  core__GEN_305_0; // @[top.scala 26:26]
  wire  core__GEN_112; // @[top.scala 26:26]
  wire  core__GEN_211; // @[top.scala 26:26]
  wire  core__GEN_220; // @[top.scala 26:26]
  wire  core__GEN_8; // @[top.scala 26:26]
  wire  core__GEN_2; // @[top.scala 26:26]
  wire  core__GEN_311_0; // @[top.scala 26:26]
  wire  core__GEN_133; // @[top.scala 26:26]
  wire  core__GEN_127; // @[top.scala 26:26]
  wire  core__GEN_288_0; // @[top.scala 26:26]
  wire  core__GEN_389; // @[top.scala 26:26]
  wire  core__GEN_91; // @[top.scala 26:26]
  wire  core__GEN_205; // @[top.scala 26:26]
  wire  core__GEN_100; // @[top.scala 26:26]
  wire  core__GEN_304; // @[top.scala 26:26]
  wire  core__GEN_60; // @[top.scala 26:26]
  wire  core__GEN_298; // @[top.scala 26:26]
  wire  core__GEN_189; // @[top.scala 26:26]
  wire  core__GEN_199; // @[top.scala 26:26]
  wire  core__GEN_177; // @[top.scala 26:26]
  wire  core__GEN_12_1; // @[top.scala 26:26]
  wire  core__GEN_268_0; // @[top.scala 26:26]
  wire  core__GEN_94; // @[top.scala 26:26]
  wire  core__GEN_376; // @[top.scala 26:26]
  wire  core__GEN_162; // @[top.scala 26:26]
  wire  core__GEN_193; // @[top.scala 26:26]
  wire  core__GEN_208; // @[top.scala 26:26]
  wire  core__GEN_454; // @[top.scala 26:26]
  wire  core__GEN_293_0; // @[top.scala 26:26]
  wire  core__GEN_261; // @[top.scala 26:26]
  wire  core__GEN_115; // @[top.scala 26:26]
  wire  core__GEN_27; // @[top.scala 26:26]
  wire  core__GEN_270; // @[top.scala 26:26]
  wire  core__GEN_392; // @[top.scala 26:26]
  wire  core__GEN_361; // @[top.scala 26:26]
  wire  core__GEN_287; // @[top.scala 26:26]
  wire  core__GEN_183; // @[top.scala 26:26]
  wire  core__GEN_256_0; // @[top.scala 26:26]
  wire  core__GEN_460; // @[top.scala 26:26]
  wire  core__GEN_278; // @[top.scala 26:26]
  wire  core__GEN_33; // @[top.scala 26:26]
  wire  core__GEN_276; // @[top.scala 26:26]
  wire  core__GEN_282_0; // @[top.scala 26:26]
  wire  core__GEN_292; // @[top.scala 26:26]
  wire  core__GEN_355; // @[top.scala 26:26]
  wire  core__GEN_48; // @[top.scala 26:26]
  wire  core__GEN_386; // @[top.scala 26:26]
  wire  core__GEN_6_1; // @[top.scala 26:26]
  wire  core__GEN_277_0; // @[top.scala 26:26]
  wire  core__GEN_21; // @[top.scala 26:26]
  wire  core__GEN_307; // @[top.scala 26:26]
  wire  core__GEN_262_0; // @[top.scala 26:26]
  wire  core__GEN_109; // @[top.scala 26:26]
  wire  core__GEN_11; // @[top.scala 26:26]
  wire  core__GEN_244_0; // @[top.scala 26:26]
  wire  core__GEN_448; // @[top.scala 26:26]
  wire  core__GEN_442; // @[top.scala 26:26]
  wire  core__GEN_21_0; // @[top.scala 26:26]
  wire  core__GEN_15_2; // @[top.scala 26:26]
  wire  core__GEN_457; // @[top.scala 26:26]
  wire  core__GEN_337; // @[top.scala 26:26]
  wire  core__GEN_30; // @[top.scala 26:26]
  wire  core__GEN_83; // @[top.scala 26:26]
  wire  core__GEN_364; // @[top.scala 26:26]
  wire  core__GEN_171; // @[top.scala 26:26]
  wire  core__GEN_186; // @[top.scala 26:26]
  wire  core__GEN_328; // @[top.scala 26:26]
  wire  core__GEN_463; // @[top.scala 26:26]
  wire  core__GEN_144; // @[top.scala 26:26]
  wire  core__GEN_279_0; // @[top.scala 26:26]
  wire  core__GEN_436; // @[top.scala 26:26]
  wire  core__GEN_97; // @[top.scala 26:26]
  wire  core__GEN_9_1; // @[top.scala 26:26]
  wire  core__GEN_264; // @[top.scala 26:26]
  wire  core__GEN_165; // @[top.scala 26:26]
  wire  core__GEN_159; // @[top.scala 26:26]
  wire  core__GEN_370; // @[top.scala 26:26]
  wire  core__GEN_250_0; // @[top.scala 26:26]
  wire  core__GEN_265_0; // @[top.scala 26:26]
  wire  core__GEN_258; // @[top.scala 26:26]
  wire  core__GEN_5; // @[top.scala 26:26]
  wire  core__GEN_285_0; // @[top.scala 26:26]
  wire  core__GEN_180; // @[top.scala 26:26]
  wire  core__GEN_271_0; // @[top.scala 26:26]
  wire  core__GEN_9_2; // @[top.scala 26:26]
  wire  core__GEN_243; // @[top.scala 26:26]
  wire  core__GEN_349; // @[top.scala 26:26]
  wire  core__GEN_343; // @[top.scala 26:26]
  wire  core__GEN_147; // @[top.scala 26:26]
  wire  core__GEN_77; // @[top.scala 26:26]
  wire  core__GEN_352; // @[top.scala 26:26]
  wire  core__GEN_174; // @[top.scala 26:26]
  wire  core__GEN_225; // @[top.scala 26:26]
  wire  core__GEN_247_0; // @[top.scala 26:26]
  wire  core__GEN_252; // @[top.scala 26:26]
  wire  core__GEN_325; // @[top.scala 26:26]
  wire  core__GEN_132; // @[top.scala 26:26]
  wire  core__GEN_147_0; // @[top.scala 26:26]
  wire  core__GEN_151_0; // @[top.scala 26:26]
  wire  core__GEN_238_0; // @[top.scala 26:26]
  wire  core__GEN_240; // @[top.scala 26:26]
  wire  core__GEN_451; // @[top.scala 26:26]
  wire  core__GEN_65; // @[top.scala 26:26]
  wire  core__GEN_273; // @[top.scala 26:26]
  wire  core__GEN_346; // @[top.scala 26:26]
  wire  core__GEN_59; // @[top.scala 26:26]
  wire  core__GEN_409; // @[top.scala 26:26]
  wire  core__GEN_231; // @[top.scala 26:26]
  wire  core__GEN_253_0; // @[top.scala 26:26]
  wire  core__GEN_331; // @[top.scala 26:26]
  wire  core__GEN_86; // @[top.scala 26:26]
  wire  core__GEN_8_0; // @[top.scala 26:26]
  wire  core__GEN_80; // @[top.scala 26:26]
  wire  core__GEN_11_0; // @[top.scala 26:26]
  wire  core__GEN_430; // @[top.scala 26:26]
  wire  core__GEN_424; // @[top.scala 26:26]
  wire  core__GEN_3_1; // @[top.scala 26:26]
  wire  core__GEN_246; // @[top.scala 26:26]
  wire  core__GEN_12_2; // @[top.scala 26:26]
  wire  core__GEN_71; // @[top.scala 26:26]
  wire  core__GEN_153; // @[top.scala 26:26]
  wire  core__GEN_168; // @[top.scala 26:26]
  wire  core__GEN_445; // @[top.scala 26:26]
  wire  core__GEN_310_0; // @[top.scala 26:26]
  wire  core__GEN_259_0; // @[top.scala 26:26]
  wire  core__GEN_267; // @[top.scala 26:26]
  wire  core__GEN_126; // @[top.scala 26:26]
  wire  core__GEN_358; // @[top.scala 26:26]
  wire  core__GEN_213; // @[top.scala 26:26]
  wire  core__GEN_255; // @[top.scala 26:26]
  wire  core__GEN_334; // @[top.scala 26:26]
  wire  core__GEN_156; // @[top.scala 26:26]
  wire  core__GEN_150; // @[top.scala 26:26]
  wire  core__GEN_412; // @[top.scala 26:26]
  wire  core__GEN_114; // @[top.scala 26:26]
  wire  core__GEN_228; // @[top.scala 26:26]
  wire  core__GEN_141; // @[top.scala 26:26]
  wire  core__GEN_11_1; // @[top.scala 26:26]
  wire  core__GEN_418; // @[top.scala 26:26]
  wire  core__GEN_427; // @[top.scala 26:26]
  wire  core__GEN_313_0; // @[top.scala 26:26]
  wire  core__GEN_292_0; // @[top.scala 26:26]
  wire  core__GEN_241_0; // @[top.scala 26:26]
  wire  core__GEN_108; // @[top.scala 26:26]
  wire  core__GEN_249; // @[top.scala 26:26]
  wire  core__GEN_6_2; // @[top.scala 26:26]
  wire  core__GEN_340; // @[top.scala 26:26]
  wire  core__GEN_312_0; // @[top.scala 26:26]
  wire  core__GEN_68; // @[top.scala 26:26]
  wire  core__GEN_74; // @[top.scala 26:26]
  wire  core__GEN_207; // @[top.scala 26:26]
  wire  core__GEN_235_0; // @[top.scala 26:26]
  wire  core__GEN_439; // @[top.scala 26:26]
  wire  core__GEN_20; // @[top.scala 26:26]
  wire  core__GEN_298_0; // @[top.scala 26:26]
  wire  core__GEN_307_0; // @[top.scala 26:26]
  wire  core__GEN_234; // @[top.scala 26:26]
  wire  core__GEN_306_0; // @[top.scala 26:26]
  wire  core__GEN_129; // @[top.scala 26:26]
  wire  core__GEN_17; // @[top.scala 26:26]
  wire  core__GEN_406; // @[top.scala 26:26]
  wire  core__GEN_89; // @[top.scala 26:26]
  wire  core__GEN_433; // @[top.scala 26:26]
  wire  core__GEN_319_0; // @[top.scala 26:26]
  wire  core__GEN_47; // @[top.scala 26:26]
  wire  core__GEN_53; // @[top.scala 26:26]
  wire  core__GEN_135; // @[top.scala 26:26]
  wire  core__GEN_391; // @[top.scala 26:26]
  wire  core__GEN_400; // @[top.scala 26:26]
  wire  core__GEN_415; // @[top.scala 26:26]
  wire  core__GEN_222; // @[top.scala 26:26]
  wire  core__GEN_295_0; // @[top.scala 26:26]
  wire  core__GEN_270_0; // @[top.scala 26:26]
  wire  core__GEN_29; // @[top.scala 26:26]
  wire  core__GEN_4_1; // @[top.scala 26:26]
  wire  core__GEN_322_0; // @[top.scala 26:26]
  wire  core__GEN_41; // @[top.scala 26:26]
  wire  core__GEN_56; // @[top.scala 26:26]
  wire  core__GEN_14; // @[top.scala 26:26]
  wire  core__GEN_195; // @[top.scala 26:26]
  wire  core__GEN_421; // @[top.scala 26:26]
  wire  core__GEN_280_0; // @[top.scala 26:26]
  wire  core__GEN_237; // @[top.scala 26:26]
  wire  core__GEN_102; // @[top.scala 26:26]
  wire  core__GEN_379; // @[top.scala 26:26]
  wire  core__GEN_62; // @[top.scala 26:26]
  wire  core__GEN_394; // @[top.scala 26:26]
  wire  core__GEN_23; // @[top.scala 26:26]
  wire  core__GEN_35; // @[top.scala 26:26]
  wire  core__GEN_123; // @[top.scala 26:26]
  wire  core__GEN_117; // @[top.scala 26:26]
  wire  core__GEN_369; // @[top.scala 26:26]
  wire  core__GEN_321; // @[top.scala 26:26]
  wire  core__GEN_216; // @[top.scala 26:26]
  wire  core__GEN_5_1; // @[top.scala 26:26]
  wire  core__GEN_14_0; // @[top.scala 26:26]
  wire  core__GEN_13_1; // @[top.scala 26:26]
  wire  core__GEN_316_0; // @[top.scala 26:26]
  wire  core__GEN_294_0; // @[top.scala 26:26]
  wire  core__GEN_50; // @[top.scala 26:26]
  wire  core__GEN_138; // @[top.scala 26:26]
  wire  core__GEN_201; // @[top.scala 26:26]
  wire  core__GEN_210; // @[top.scala 26:26]
  wire  core__GEN_96; // @[top.scala 26:26]
  wire  core__GEN_301_0; // @[top.scala 26:26]
  wire  core__GEN_315; // @[top.scala 26:26]
  wire  core__GEN_309; // @[top.scala 26:26]
  wire  core__GEN_17_0; // @[top.scala 26:26]
  wire  core__GEN_283_0; // @[top.scala 26:26]
  wire  core__GEN_273_0; // @[top.scala 26:26]
  wire  core__GEN_105; // @[top.scala 26:26]
  wire  core__GEN_382; // @[top.scala 26:26]
  wire  core__GEN_303; // @[top.scala 26:26]
  wire  core__GEN_204; // @[top.scala 26:26]
  wire  core__GEN_318_0; // @[top.scala 26:26]
  wire  core__GEN_173; // @[top.scala 26:26]
  wire  core__GEN_198; // @[top.scala 26:26]
  wire  core__GEN_258_0; // @[top.scala 26:26]
  wire  core__GEN_304_0; // @[top.scala 26:26]
  wire  core__GEN_23_0; // @[top.scala 26:26]
  wire  core__GEN_272_0; // @[top.scala 26:26]
  wire  core__GEN_120; // @[top.scala 26:26]
  wire  core__GEN_403; // @[top.scala 26:26]
  wire  core__GEN_372; // @[top.scala 26:26]
  wire  core__GEN_366; // @[top.scala 26:26]
  wire  core__GEN_267_0; // @[top.scala 26:26]
  wire  core__GEN_188; // @[top.scala 26:26]
  wire  core__GEN_289_0; // @[top.scala 26:26]
  wire  core__GEN_1_2; // @[top.scala 26:26]
  wire  core__GEN_44; // @[top.scala 26:26]
  wire  core__GEN_287_0; // @[top.scala 26:26]
  wire  core__GEN_297; // @[top.scala 26:26]
  wire  core__GEN_388; // @[top.scala 26:26]
  wire  core__GEN_397; // @[top.scala 26:26]
  wire  core__GEN_2_1; // @[top.scala 26:26]
  wire  core__GEN_252_0; // @[top.scala 26:26]
  wire  core__GEN_450; // @[top.scala 26:26]
  wire  core__GEN_99; // @[top.scala 26:26]
  wire  core__GEN_351; // @[top.scala 26:26]
  wire  core__GEN_38; // @[top.scala 26:26]
  wire  core__GEN_111; // @[top.scala 26:26]
  wire  core__GEN_219; // @[top.scala 26:26]
  wire  core__GEN_17_1; // @[top.scala 26:26]
  wire  core__GEN_7_1; // @[top.scala 26:26]
  wire  core__GEN_453; // @[top.scala 26:26]
  wire  core__GEN_447; // @[top.scala 26:26]
  wire  core__GEN_26; // @[top.scala 26:26]
  wire  core__GEN_176; // @[top.scala 26:26]
  wire  core__GEN_182; // @[top.scala 26:26]
  wire  core__GEN_438; // @[top.scala 26:26]
  wire  core__GEN_333; // @[top.scala 26:26]
  wire  core__GEN_290_0; // @[top.scala 26:26]
  wire  core__GEN_240_0; // @[top.scala 26:26]
  wire  core__GEN_0_1; // @[top.scala 26:26]
  wire  core__GEN_339; // @[top.scala 26:26]
  wire  core__GEN_32; // @[top.scala 26:26]
  wire  core__GEN_161; // @[top.scala 26:26]
  wire  core__GEN_275_0; // @[top.scala 26:26]
  wire  core__GEN_170; // @[top.scala 26:26]
  wire  core__GEN_375; // @[top.scala 26:26]
  wire  core__GEN_261_0; // @[top.scala 26:26]
  wire  core__GEN_192; // @[top.scala 26:26]
  wire  core__GEN_20_0; // @[top.scala 26:26]
  wire  core__GEN_255_0; // @[top.scala 26:26]
  wire  core__GEN_269_0; // @[top.scala 26:26]
  wire  core__GEN_10_2; // @[top.scala 26:26]
  wire  core__GEN_360; // @[top.scala 26:26]
  wire  core__GEN_281_0; // @[top.scala 26:26]
  wire  core__GEN_291_0; // @[top.scala 26:26]
  wire  core__GEN_155; // @[top.scala 26:26]
  wire  core__GEN_88; // @[top.scala 26:26]
  wire  core__GEN_300_0; // @[top.scala 26:26]
  wire  core__GEN_432; // @[top.scala 26:26]
  wire  core__GEN_11_2; // @[top.scala 26:26]
  wire  core__GEN_286_0; // @[top.scala 26:26]
  wire  core__GEN_276_0; // @[top.scala 26:26]
  wire  core__GEN_5_2; // @[top.scala 26:26]
  wire  core__GEN_254_0; // @[top.scala 26:26]
  wire  core__GEN_93; // @[top.scala 26:26]
  wire  core__GEN_5_3; // @[top.scala 26:26]
  wire  core__GEN_459; // @[top.scala 26:26]
  wire  core__GEN_385; // @[top.scala 26:26]
  wire  core__GEN_354; // @[top.scala 26:26]
  wire  core__GEN_234_0; // @[top.scala 26:26]
  wire  core__GEN_3_2; // @[top.scala 26:26]
  wire  core__GEN_146; // @[top.scala 26:26]
  wire  core__GEN_441; // @[top.scala 26:26]
  wire  core__GEN_321_0; // @[top.scala 26:26]
  wire  core__GEN_14_1; // @[top.scala 26:26]
  wire  core__GEN_257_0; // @[top.scala 26:26]
  wire  core__GEN_13_2; // @[top.scala 26:26]
  wire  core__GEN_348; // @[top.scala 26:26]
  wire  core__GEN_82; // @[top.scala 26:26]
  wire  core__GEN_357; // @[top.scala 26:26]
  wire  core__GEN_243_0; // @[top.scala 26:26]
  wire  core__GEN_8_1; // @[top.scala 26:26]
  wire  core__GEN_8_2; // @[top.scala 26:26]
  wire  core__GEN_462; // @[top.scala 26:26]
  wire  core__GEN_456; // @[top.scala 26:26]
  wire  core__GEN_342; // @[top.scala 26:26]
  wire  core__GEN_278_0; // @[top.scala 26:26]
  wire  core__GEN_70; // @[top.scala 26:26]
  wire  core__GEN_158; // @[top.scala 26:26]
  wire  core__GEN_420; // @[top.scala 26:26]
  wire  core__GEN_414; // @[top.scala 26:26]
  wire  core__GEN_236_0; // @[top.scala 26:26]
  wire  core__GEN_185; // @[top.scala 26:26]
  wire  core__GEN_336; // @[top.scala 26:26]
  wire  core__GEN_61; // @[top.scala 26:26]
  wire  core__GEN_143; // @[top.scala 26:26]
  wire  core__GEN_284_0; // @[top.scala 26:26]
  wire  core__GEN_179; // @[top.scala 26:26]
  wire  core__GEN_435; // @[top.scala 26:26]
  wire  core__GEN_242_0; // @[top.scala 26:26]
  wire  core__GEN_249_0; // @[top.scala 26:26]
  wire  core__GEN_137; // @[top.scala 26:26]
  wire  core__GEN_76; // @[top.scala 26:26]
  wire  core__GEN_164; // @[top.scala 26:26]
  wire  core__GEN_237_0; // @[top.scala 26:26]
  wire  core__GEN_315_0; // @[top.scala 26:26]
  wire  core__GEN_264_0; // @[top.scala 26:26]
  wire  core__GEN_263_0; // @[top.scala 26:26]
  wire  core__GEN_363; // @[top.scala 26:26]
  wire  core__GEN_167; // @[top.scala 26:26]
  wire  core__GEN_246_0; // @[top.scala 26:26]
  wire  core__GEN_43; // @[top.scala 26:26]
  wire  core__GEN_266_0; // @[top.scala 26:26]
  wire  core__GEN_131; // @[top.scala 26:26]
  wire  core__GEN_125; // @[top.scala 26:26]
  wire  core__GEN_317_0; // @[top.scala 26:26]
  wire  core__GEN_224; // @[top.scala 26:26]
  wire  core__GEN_150_0; // @[top.scala 26:26]
  wire  core__GEN_119; // @[top.scala 26:26]
  wire  core__GEN_239_0; // @[top.scala 26:26]
  wire  core__GEN_330; // @[top.scala 26:26]
  wire  core__GEN_152_0; // @[top.scala 26:26]
  wire  core__GEN_146_0; // @[top.scala 26:26]
  wire  core__GEN_7_2; // @[top.scala 26:26]
  wire  core__GEN_297_0; // @[top.scala 26:26]
  wire  core__GEN_245_0; // @[top.scala 26:26]
  wire  core__GEN_11_3; // @[top.scala 26:26]
  wire  core__GEN_345; // @[top.scala 26:26]
  wire  core__GEN_323_0; // @[top.scala 26:26]
  wire  core__GEN_396; // @[top.scala 26:26]
  wire  core__GEN_79; // @[top.scala 26:26]
  wire  core__GEN_218; // @[top.scala 26:26]
  wire  core__GEN_408; // @[top.scala 26:26]
  wire  core__GEN_423; // @[top.scala 26:26]
  wire  core__GEN_309_0; // @[top.scala 26:26]
  wire  core__GEN_303_0; // @[top.scala 26:26]
  wire  core__GEN_64; // @[top.scala 26:26]
  wire  core__GEN_417; // @[top.scala 26:26]
  wire  core__GEN_429; // @[top.scala 26:26]
  wire  core__GEN_444; // @[top.scala 26:26]
  wire  core__GEN_324; // @[top.scala 26:26]
  wire  core__GEN_58; // @[top.scala 26:26]
  wire  core__GEN_251_0; // @[top.scala 26:26]
  wire  core__GEN_260_0; // @[top.scala 26:26]
  wire  core__GEN_140; // @[top.scala 26:26]
  wire  core__GEN_402; // @[top.scala 26:26]
  wire  core__GEN_85; // @[top.scala 26:26]
  wire  memory_metaReset; // @[top.scala 29:28]
  wire  memory_clock; // @[top.scala 29:28]
  wire [31:0] memory_io_core_ports_0_req_bits_addr; // @[top.scala 29:28]
  wire [31:0] memory_io_core_ports_0_req_bits_data; // @[top.scala 29:28]
  wire  memory_io_core_ports_0_req_bits_fcn; // @[top.scala 29:28]
  wire [2:0] memory_io_core_ports_0_req_bits_typ; // @[top.scala 29:28]
  wire [31:0] memory_io_core_ports_0_resp_bits_data; // @[top.scala 29:28]
  wire  memory__GEN_1_0; // @[top.scala 29:28]
  wire  memory__GEN_4_0; // @[top.scala 29:28]
  wire  memory__GEN_0_1; // @[top.scala 29:28]
  wire  memory__GEN_3_1; // @[top.scala 29:28]
  wire  memory__GEN_2_1; // @[top.scala 29:28]
  wire  memory__GEN_5_1; // @[top.scala 29:28]
  wire  profilePin = core__GEN_1_0;
  wire  profilePin_0 = core__GEN_5_3;
  wire  profilePin_1 = core__GEN_6_2;
  wire  profilePin_2 = core__GEN_7_0;
  wire  profilePin_3 = core__GEN_8_2;
  wire  profilePin_4 = core__GEN_9_1;
  wire  profilePin_5 = core__GEN_10_0;
  wire  profilePin_6 = core__GEN_11_3;
  wire  profilePin_7 = core__GEN_12_2;
  wire  profilePin_8 = core__GEN_13_0;
  wire [9:0] _GEN_627 = {profilePin,profilePin_0,profilePin_1,profilePin_2,profilePin_3,profilePin_4,profilePin_5,profilePin_6,profilePin_7,profilePin_8};
  wire  profilePin_9 = core__GEN_0_1;
  wire  profilePin_10 = core__GEN_1_1;
  wire  profilePin_11 = core__GEN_2_1;
  wire  profilePin_12 = core__GEN_3_1;
  wire  profilePin_13 = core__GEN_4_0;
  wire  profilePin_14 = core__GEN_5_2;
  wire  profilePin_15 = core__GEN_6_1;
  wire  profilePin_16 = core__GEN_7;
  wire  profilePin_17 = core__GEN_8_1;
  wire [18:0] _GEN_636 = {_GEN_627,profilePin_9,profilePin_10,profilePin_11,profilePin_12,profilePin_13,profilePin_14,profilePin_15,profilePin_16,profilePin_17};
  wire  profilePin_18 = core__GEN_9_2;
  wire  profilePin_19 = core__GEN_10_1;
  wire  profilePin_20 = core__GEN_11_2;
  wire  profilePin_21 = core__GEN_12_1;
  wire  profilePin_22 = core__GEN_13;
  wire  profilePin_23 = core__GEN_14_1;
  wire  profilePin_24 = core__GEN_15_2;
  wire  profilePin_25 = core__GEN_16_1;
  wire  profilePin_26 = core__GEN_17_0;
  wire [27:0] _GEN_645 = {_GEN_636,profilePin_18,profilePin_19,profilePin_20,profilePin_21,profilePin_22,profilePin_23,profilePin_24,profilePin_25,profilePin_26};
  wire  profilePin_27 = core__GEN_18_0;
  wire  profilePin_28 = core__GEN_19_0;
  wire  profilePin_29 = core__GEN_20_0;
  wire  profilePin_30 = core__GEN_21_0;
  wire  profilePin_31 = core__GEN_22_0;
  wire  profilePin_32 = core__GEN_23_0;
  wire  profilePin_33 = core__GEN_24;
  wire  profilePin_34 = core__GEN_25;
  wire  profilePin_35 = core__GEN_26;
  wire [36:0] _GEN_654 = {_GEN_645,profilePin_27,profilePin_28,profilePin_29,profilePin_30,profilePin_31,profilePin_32,profilePin_33,profilePin_34,profilePin_35};
  wire  profilePin_36 = core__GEN_27;
  wire  profilePin_37 = core__GEN_28;
  wire  profilePin_38 = core__GEN_29;
  wire  profilePin_39 = core__GEN_30;
  wire  profilePin_40 = core__GEN_31;
  wire  profilePin_41 = core__GEN_32;
  wire  profilePin_42 = core__GEN_33;
  wire  profilePin_43 = core__GEN_34;
  wire  profilePin_44 = core__GEN_35;
  wire [45:0] _GEN_663 = {_GEN_654,profilePin_36,profilePin_37,profilePin_38,profilePin_39,profilePin_40,profilePin_41,profilePin_42,profilePin_43,profilePin_44};
  wire  profilePin_45 = core__GEN_36;
  wire  profilePin_46 = core__GEN_37;
  wire  profilePin_47 = core__GEN_38;
  wire  profilePin_48 = core__GEN_39;
  wire  profilePin_49 = core__GEN_40;
  wire  profilePin_50 = core__GEN_41;
  wire  profilePin_51 = core__GEN_42;
  wire  profilePin_52 = core__GEN_43;
  wire  profilePin_53 = core__GEN_44;
  wire [54:0] _GEN_672 = {_GEN_663,profilePin_45,profilePin_46,profilePin_47,profilePin_48,profilePin_49,profilePin_50,profilePin_51,profilePin_52,profilePin_53};
  wire  profilePin_54 = core__GEN_45;
  wire  profilePin_55 = core__GEN_46;
  wire  profilePin_56 = core__GEN_47;
  wire  profilePin_57 = core__GEN_48;
  wire  profilePin_58 = core__GEN_49;
  wire  profilePin_59 = core__GEN_50;
  wire  profilePin_60 = core__GEN_51;
  wire  profilePin_61 = core__GEN_52;
  wire  profilePin_62 = core__GEN_53;
  wire [63:0] _GEN_681 = {_GEN_672,profilePin_54,profilePin_55,profilePin_56,profilePin_57,profilePin_58,profilePin_59,profilePin_60,profilePin_61,profilePin_62};
  wire  profilePin_63 = core__GEN_54;
  wire  profilePin_64 = core__GEN_55;
  wire  profilePin_65 = core__GEN_56;
  wire  profilePin_66 = core__GEN_57;
  wire  profilePin_67 = core__GEN_58;
  wire  profilePin_68 = core__GEN_59;
  wire  profilePin_69 = core__GEN_60;
  wire  profilePin_70 = core__GEN_61;
  wire  profilePin_71 = core__GEN_62;
  wire [72:0] _GEN_690 = {_GEN_681,profilePin_63,profilePin_64,profilePin_65,profilePin_66,profilePin_67,profilePin_68,profilePin_69,profilePin_70,profilePin_71};
  wire  profilePin_72 = core__GEN_63;
  wire  profilePin_73 = core__GEN_64;
  wire  profilePin_74 = core__GEN_65;
  wire  profilePin_75 = core__GEN_66;
  wire  profilePin_76 = core__GEN_67;
  wire  profilePin_77 = core__GEN_68;
  wire  profilePin_78 = core__GEN_69;
  wire  profilePin_79 = core__GEN_70;
  wire  profilePin_80 = core__GEN_71;
  wire [81:0] _GEN_699 = {_GEN_690,profilePin_72,profilePin_73,profilePin_74,profilePin_75,profilePin_76,profilePin_77,profilePin_78,profilePin_79,profilePin_80};
  wire  profilePin_81 = core__GEN_72;
  wire  profilePin_82 = core__GEN_73;
  wire  profilePin_83 = core__GEN_74;
  wire  profilePin_84 = core__GEN_75;
  wire  profilePin_85 = core__GEN_76;
  wire  profilePin_86 = core__GEN_77;
  wire  profilePin_87 = core__GEN_78;
  wire  profilePin_88 = core__GEN_79;
  wire  profilePin_89 = core__GEN_80;
  wire [90:0] _GEN_708 = {_GEN_699,profilePin_81,profilePin_82,profilePin_83,profilePin_84,profilePin_85,profilePin_86,profilePin_87,profilePin_88,profilePin_89};
  wire  profilePin_90 = core__GEN_81;
  wire  profilePin_91 = core__GEN_82;
  wire  profilePin_92 = core__GEN_83;
  wire  profilePin_93 = core__GEN_84;
  wire  profilePin_94 = core__GEN_85;
  wire  profilePin_95 = core__GEN_86;
  wire  profilePin_96 = core__GEN_87;
  wire  profilePin_97 = core__GEN_88;
  wire  profilePin_98 = core__GEN_89;
  wire [99:0] _GEN_717 = {_GEN_708,profilePin_90,profilePin_91,profilePin_92,profilePin_93,profilePin_94,profilePin_95,profilePin_96,profilePin_97,profilePin_98};
  wire  profilePin_99 = core__GEN_90;
  wire  profilePin_100 = core__GEN_91;
  wire  profilePin_101 = core__GEN_92;
  wire  profilePin_102 = core__GEN_93;
  wire  profilePin_103 = core__GEN_94;
  wire  profilePin_104 = core__GEN_95;
  wire  profilePin_105 = core__GEN_96;
  wire  profilePin_106 = core__GEN_97;
  wire  profilePin_107 = core__GEN_98;
  wire [108:0] _GEN_726 = {_GEN_717,profilePin_99,profilePin_100,profilePin_101,profilePin_102,profilePin_103,profilePin_104,profilePin_105,profilePin_106,profilePin_107};
  wire  profilePin_108 = core__GEN_99;
  wire  profilePin_109 = core__GEN_100;
  wire  profilePin_110 = core__GEN_101;
  wire  profilePin_111 = core__GEN_102;
  wire  profilePin_112 = core__GEN_103;
  wire  profilePin_113 = core__GEN_104;
  wire  profilePin_114 = core__GEN_105;
  wire  profilePin_115 = core__GEN_106;
  wire  profilePin_116 = core__GEN_107;
  wire [117:0] _GEN_735 = {_GEN_726,profilePin_108,profilePin_109,profilePin_110,profilePin_111,profilePin_112,profilePin_113,profilePin_114,profilePin_115,profilePin_116};
  wire  profilePin_117 = core__GEN_108;
  wire  profilePin_118 = core__GEN_109;
  wire  profilePin_119 = core__GEN_110;
  wire  profilePin_120 = core__GEN_111;
  wire  profilePin_121 = core__GEN_112;
  wire  profilePin_122 = core__GEN_113;
  wire  profilePin_123 = core__GEN_114;
  wire  profilePin_124 = core__GEN_115;
  wire  profilePin_125 = core__GEN_116;
  wire [126:0] _GEN_744 = {_GEN_735,profilePin_117,profilePin_118,profilePin_119,profilePin_120,profilePin_121,profilePin_122,profilePin_123,profilePin_124,profilePin_125};
  wire  profilePin_126 = core__GEN_117;
  wire  profilePin_127 = core__GEN_118;
  wire  profilePin_128 = core__GEN_119;
  wire  profilePin_129 = core__GEN_120;
  wire  profilePin_130 = core__GEN_121;
  wire  profilePin_131 = core__GEN_122;
  wire  profilePin_132 = core__GEN_123;
  wire  profilePin_133 = core__GEN_124;
  wire  profilePin_134 = core__GEN_125;
  wire [135:0] _GEN_753 = {_GEN_744,profilePin_126,profilePin_127,profilePin_128,profilePin_129,profilePin_130,profilePin_131,profilePin_132,profilePin_133,profilePin_134};
  wire  profilePin_135 = core__GEN_126;
  wire  profilePin_136 = core__GEN_127;
  wire  profilePin_137 = core__GEN_128;
  wire  profilePin_138 = core__GEN_129;
  wire  profilePin_139 = core__GEN_130;
  wire  profilePin_140 = core__GEN_131;
  wire  profilePin_141 = core__GEN_132;
  wire  profilePin_142 = core__GEN_133;
  wire  profilePin_143 = core__GEN_134;
  wire [144:0] _GEN_762 = {_GEN_753,profilePin_135,profilePin_136,profilePin_137,profilePin_138,profilePin_139,profilePin_140,profilePin_141,profilePin_142,profilePin_143};
  wire  profilePin_144 = core__GEN_135;
  wire  profilePin_145 = core__GEN_136;
  wire  profilePin_146 = core__GEN_137;
  wire  profilePin_147 = core__GEN_138;
  wire  profilePin_148 = core__GEN_139;
  wire  profilePin_149 = core__GEN_140;
  wire  profilePin_150 = core__GEN_141;
  wire  profilePin_151 = core__GEN_142;
  wire  profilePin_152 = core__GEN_143;
  wire [153:0] _GEN_771 = {_GEN_762,profilePin_144,profilePin_145,profilePin_146,profilePin_147,profilePin_148,profilePin_149,profilePin_150,profilePin_151,profilePin_152};
  wire  profilePin_153 = core__GEN_144;
  wire  profilePin_154 = core__GEN_145;
  wire  profilePin_155 = core__GEN_146_0;
  wire  profilePin_156 = core__GEN_147_0;
  wire  profilePin_157 = core__GEN_148;
  wire  profilePin_158 = core__GEN_149;
  wire  profilePin_159 = core__GEN_150;
  wire  profilePin_160 = core__GEN_151;
  wire  profilePin_161 = core__GEN_152_0;
  wire [162:0] _GEN_780 = {_GEN_771,profilePin_153,profilePin_154,profilePin_155,profilePin_156,profilePin_157,profilePin_158,profilePin_159,profilePin_160,profilePin_161};
  wire  profilePin_162 = core__GEN_153;
  wire  profilePin_163 = core__GEN_154;
  wire  profilePin_164 = core__GEN_155;
  wire  profilePin_165 = core__GEN_156;
  wire  profilePin_166 = core__GEN_157;
  wire  profilePin_167 = core__GEN_158;
  wire  profilePin_168 = core__GEN_159;
  wire  profilePin_169 = core__GEN_160;
  wire  profilePin_170 = core__GEN_161;
  wire [171:0] _GEN_789 = {_GEN_780,profilePin_162,profilePin_163,profilePin_164,profilePin_165,profilePin_166,profilePin_167,profilePin_168,profilePin_169,profilePin_170};
  wire  profilePin_171 = core__GEN_162;
  wire  profilePin_172 = core__GEN_163;
  wire  profilePin_173 = core__GEN_164;
  wire  profilePin_174 = core__GEN_165;
  wire  profilePin_175 = core__GEN_166;
  wire  profilePin_176 = core__GEN_167;
  wire  profilePin_177 = core__GEN_168;
  wire  profilePin_178 = core__GEN_169;
  wire  profilePin_179 = core__GEN_170;
  wire [180:0] _GEN_798 = {_GEN_789,profilePin_171,profilePin_172,profilePin_173,profilePin_174,profilePin_175,profilePin_176,profilePin_177,profilePin_178,profilePin_179};
  wire  profilePin_180 = core__GEN_171;
  wire  profilePin_181 = core__GEN_172;
  wire  profilePin_182 = core__GEN_173;
  wire  profilePin_183 = core__GEN_174;
  wire  profilePin_184 = core__GEN_175;
  wire  profilePin_185 = core__GEN_176;
  wire  profilePin_186 = core__GEN_177;
  wire  profilePin_187 = core__GEN_178;
  wire  profilePin_188 = core__GEN_179;
  wire [189:0] _GEN_807 = {_GEN_798,profilePin_180,profilePin_181,profilePin_182,profilePin_183,profilePin_184,profilePin_185,profilePin_186,profilePin_187,profilePin_188};
  wire  profilePin_189 = core__GEN_180;
  wire  profilePin_190 = core__GEN_181;
  wire  profilePin_191 = core__GEN_182;
  wire  profilePin_192 = core__GEN_183;
  wire  profilePin_193 = core__GEN_184;
  wire  profilePin_194 = core__GEN_185;
  wire  profilePin_195 = core__GEN_186;
  wire  profilePin_196 = core__GEN_187;
  wire  profilePin_197 = core__GEN_188;
  wire [198:0] _GEN_816 = {_GEN_807,profilePin_189,profilePin_190,profilePin_191,profilePin_192,profilePin_193,profilePin_194,profilePin_195,profilePin_196,profilePin_197};
  wire  profilePin_198 = core__GEN_189;
  wire  profilePin_199 = core__GEN_190;
  wire  profilePin_200 = core__GEN_191;
  wire  profilePin_201 = core__GEN_192;
  wire  profilePin_202 = core__GEN_193;
  wire  profilePin_203 = core__GEN_194;
  wire  profilePin_204 = core__GEN_195;
  wire  profilePin_205 = core__GEN_196;
  wire  profilePin_206 = core__GEN_197;
  wire [207:0] _GEN_825 = {_GEN_816,profilePin_198,profilePin_199,profilePin_200,profilePin_201,profilePin_202,profilePin_203,profilePin_204,profilePin_205,profilePin_206};
  wire  profilePin_207 = core__GEN_198;
  wire  profilePin_208 = core__GEN_199;
  wire  profilePin_209 = core__GEN_200;
  wire  profilePin_210 = core__GEN_201;
  wire  profilePin_211 = core__GEN_202;
  wire  profilePin_212 = core__GEN_203;
  wire  profilePin_213 = core__GEN_204;
  wire  profilePin_214 = core__GEN_205;
  wire  profilePin_215 = core__GEN_206;
  wire [216:0] _GEN_834 = {_GEN_825,profilePin_207,profilePin_208,profilePin_209,profilePin_210,profilePin_211,profilePin_212,profilePin_213,profilePin_214,profilePin_215};
  wire  profilePin_216 = core__GEN_207;
  wire  profilePin_217 = core__GEN_208;
  wire  profilePin_218 = core__GEN_209;
  wire  profilePin_219 = core__GEN_210;
  wire  profilePin_220 = core__GEN_211;
  wire  profilePin_221 = core__GEN_212;
  wire  profilePin_222 = core__GEN_213;
  wire  profilePin_223 = core__GEN_214;
  wire  profilePin_224 = core__GEN_215;
  wire [225:0] _GEN_843 = {_GEN_834,profilePin_216,profilePin_217,profilePin_218,profilePin_219,profilePin_220,profilePin_221,profilePin_222,profilePin_223,profilePin_224};
  wire  profilePin_225 = core__GEN_216;
  wire  profilePin_226 = core__GEN_217;
  wire  profilePin_227 = core__GEN_218;
  wire  profilePin_228 = core__GEN_219;
  wire  profilePin_229 = core__GEN_220;
  wire  profilePin_230 = core__GEN_221;
  wire  profilePin_231 = core__GEN_222;
  wire  profilePin_232 = core__GEN_223;
  wire  profilePin_233 = core__GEN_224;
  wire [234:0] _GEN_852 = {_GEN_843,profilePin_225,profilePin_226,profilePin_227,profilePin_228,profilePin_229,profilePin_230,profilePin_231,profilePin_232,profilePin_233};
  wire  profilePin_234 = core__GEN_225;
  wire  profilePin_235 = core__GEN_226;
  wire  profilePin_236 = core__GEN_227;
  wire  profilePin_237 = core__GEN_228;
  wire  profilePin_238 = core__GEN_229;
  wire  profilePin_239 = core__GEN_230;
  wire  profilePin_240 = core__GEN_231;
  wire  profilePin_241 = core__GEN_232;
  wire  profilePin_242 = core__GEN_233;
  wire [243:0] _GEN_861 = {_GEN_852,profilePin_234,profilePin_235,profilePin_236,profilePin_237,profilePin_238,profilePin_239,profilePin_240,profilePin_241,profilePin_242};
  wire  profilePin_243 = core__GEN_234;
  wire  profilePin_244 = core__GEN_235;
  wire  profilePin_245 = core__GEN_236_0;
  wire  profilePin_246 = core__GEN_237;
  wire  profilePin_247 = core__GEN_238;
  wire  profilePin_248 = core__GEN_239_0;
  wire  profilePin_249 = core__GEN_240;
  wire  profilePin_250 = core__GEN_241;
  wire  profilePin_251 = core__GEN_242_0;
  wire [252:0] _GEN_870 = {_GEN_861,profilePin_243,profilePin_244,profilePin_245,profilePin_246,profilePin_247,profilePin_248,profilePin_249,profilePin_250,profilePin_251};
  wire  profilePin_252 = core__GEN_243;
  wire  profilePin_253 = core__GEN_244;
  wire  profilePin_254 = core__GEN_245_0;
  wire  profilePin_255 = core__GEN_246;
  wire  profilePin_256 = core__GEN_247;
  wire  profilePin_257 = core__GEN_248;
  wire  profilePin_258 = core__GEN_249;
  wire  profilePin_259 = core__GEN_250;
  wire  profilePin_260 = core__GEN_251_0;
  wire [261:0] _GEN_879 = {_GEN_870,profilePin_252,profilePin_253,profilePin_254,profilePin_255,profilePin_256,profilePin_257,profilePin_258,profilePin_259,profilePin_260};
  wire  profilePin_261 = core__GEN_252;
  wire  profilePin_262 = core__GEN_253;
  wire  profilePin_263 = core__GEN_254_0;
  wire  profilePin_264 = core__GEN_255;
  wire  profilePin_265 = core__GEN_256;
  wire  profilePin_266 = core__GEN_257_0;
  wire  profilePin_267 = core__GEN_258;
  wire  profilePin_268 = core__GEN_259;
  wire  profilePin_269 = core__GEN_260_0;
  wire [270:0] _GEN_888 = {_GEN_879,profilePin_261,profilePin_262,profilePin_263,profilePin_264,profilePin_265,profilePin_266,profilePin_267,profilePin_268,profilePin_269};
  wire  profilePin_270 = core__GEN_261;
  wire  profilePin_271 = core__GEN_262;
  wire  profilePin_272 = core__GEN_263_0;
  wire  profilePin_273 = core__GEN_264;
  wire  profilePin_274 = core__GEN_265;
  wire  profilePin_275 = core__GEN_266_0;
  wire  profilePin_276 = core__GEN_267;
  wire  profilePin_277 = core__GEN_268;
  wire  profilePin_278 = core__GEN_269_0;
  wire [279:0] _GEN_897 = {_GEN_888,profilePin_270,profilePin_271,profilePin_272,profilePin_273,profilePin_274,profilePin_275,profilePin_276,profilePin_277,profilePin_278};
  wire  profilePin_279 = core__GEN_270;
  wire  profilePin_280 = core__GEN_271;
  wire  profilePin_281 = core__GEN_272_0;
  wire  profilePin_282 = core__GEN_273;
  wire  profilePin_283 = core__GEN_274;
  wire  profilePin_284 = core__GEN_275_0;
  wire  profilePin_285 = core__GEN_276;
  wire  profilePin_286 = core__GEN_277;
  wire  profilePin_287 = core__GEN_278_0;
  wire [288:0] _GEN_906 = {_GEN_897,profilePin_279,profilePin_280,profilePin_281,profilePin_282,profilePin_283,profilePin_284,profilePin_285,profilePin_286,profilePin_287};
  wire  profilePin_288 = core__GEN_279_0;
  wire  profilePin_289 = core__GEN_280;
  wire  profilePin_290 = core__GEN_281_0;
  wire  profilePin_291 = core__GEN_282_0;
  wire  profilePin_292 = core__GEN_283;
  wire  profilePin_293 = core__GEN_284_0;
  wire  profilePin_294 = core__GEN_285_0;
  wire  profilePin_295 = core__GEN_286;
  wire  profilePin_296 = core__GEN_287_0;
  wire [297:0] _GEN_915 = {_GEN_906,profilePin_288,profilePin_289,profilePin_290,profilePin_291,profilePin_292,profilePin_293,profilePin_294,profilePin_295,profilePin_296};
  wire  profilePin_297 = core__GEN_288_0;
  wire  profilePin_298 = core__GEN_289;
  wire  profilePin_299 = core__GEN_290_0;
  wire  profilePin_300 = core__GEN_291_0;
  wire  profilePin_301 = core__GEN_292;
  wire  profilePin_302 = core__GEN_293;
  wire  profilePin_303 = core__GEN_294_0;
  wire  profilePin_304 = core__GEN_295;
  wire  profilePin_305 = core__GEN_296;
  wire [306:0] _GEN_924 = {_GEN_915,profilePin_297,profilePin_298,profilePin_299,profilePin_300,profilePin_301,profilePin_302,profilePin_303,profilePin_304,profilePin_305};
  wire  profilePin_306 = core__GEN_297;
  wire  profilePin_307 = core__GEN_298;
  wire  profilePin_308 = core__GEN_299;
  wire  profilePin_309 = core__GEN_300_0;
  wire  profilePin_310 = core__GEN_301;
  wire  profilePin_311 = core__GEN_302;
  wire  profilePin_312 = core__GEN_303;
  wire  profilePin_313 = core__GEN_304;
  wire  profilePin_314 = core__GEN_305;
  wire [315:0] _GEN_933 = {_GEN_924,profilePin_306,profilePin_307,profilePin_308,profilePin_309,profilePin_310,profilePin_311,profilePin_312,profilePin_313,profilePin_314};
  wire  profilePin_315 = core__GEN_306_0;
  wire  profilePin_316 = core__GEN_307;
  wire  profilePin_317 = core__GEN_308;
  wire  profilePin_318 = core__GEN_309;
  wire  profilePin_319 = core__GEN_310;
  wire  profilePin_320 = core__GEN_311;
  wire  profilePin_321 = core__GEN_312_0;
  wire  profilePin_322 = core__GEN_313;
  wire  profilePin_323 = core__GEN_314;
  wire [324:0] _GEN_942 = {_GEN_933,profilePin_315,profilePin_316,profilePin_317,profilePin_318,profilePin_319,profilePin_320,profilePin_321,profilePin_322,profilePin_323};
  wire  profilePin_324 = core__GEN_315;
  wire  profilePin_325 = core__GEN_316;
  wire  profilePin_326 = core__GEN_317_0;
  wire  profilePin_327 = core__GEN_318_0;
  wire  profilePin_328 = core__GEN_319;
  wire  profilePin_329 = core__GEN_320;
  wire  profilePin_330 = core__GEN_321;
  wire  profilePin_331 = core__GEN_322;
  wire  profilePin_332 = core__GEN_323_0;
  wire [333:0] _GEN_951 = {_GEN_942,profilePin_324,profilePin_325,profilePin_326,profilePin_327,profilePin_328,profilePin_329,profilePin_330,profilePin_331,profilePin_332};
  wire  profilePin_333 = core__GEN_8_0;
  wire  profilePin_334 = core__GEN_9_0;
  wire  profilePin_335 = core__GEN_10;
  wire  profilePin_336 = core__GEN_11_1;
  wire  profilePin_337 = core__GEN_12_0;
  wire  profilePin_338 = core__GEN_13_2;
  wire  profilePin_339 = core__GEN_14;
  wire  profilePin_340 = core__GEN_15_0;
  wire  profilePin_341 = core__GEN_16;
  wire [342:0] _GEN_960 = {_GEN_951,profilePin_333,profilePin_334,profilePin_335,profilePin_336,profilePin_337,profilePin_338,profilePin_339,profilePin_340,profilePin_341};
  wire  profilePin_342 = core__GEN_17;
  wire  profilePin_343 = core__GEN_18;
  wire  profilePin_344 = core__GEN_3_2;
  wire  profilePin_345 = core__GEN_5_1;
  wire  profilePin_346 = core__GEN_6_0;
  wire  profilePin_347 = core__GEN_7_2;
  wire  profilePin_348 = core__GEN_11_0;
  wire  profilePin_349 = core__GEN_15;
  wire  profilePin_350 = core__GEN_146;
  wire [351:0] _GEN_969 = {_GEN_960,profilePin_342,profilePin_343,profilePin_344,profilePin_345,profilePin_346,profilePin_347,profilePin_348,profilePin_349,profilePin_350};
  wire  profilePin_351 = core__GEN_147;
  wire  profilePin_352 = core__GEN_149_0;
  wire  profilePin_353 = core__GEN_150_0;
  wire  profilePin_354 = core__GEN_151_0;
  wire  profilePin_355 = core__GEN_152;
  wire  profilePin_356 = core__GEN_234_0;
  wire  profilePin_357 = core__GEN_235_0;
  wire  profilePin_358 = core__GEN_236;
  wire  profilePin_359 = core__GEN_237_0;
  wire [360:0] _GEN_978 = {_GEN_969,profilePin_351,profilePin_352,profilePin_353,profilePin_354,profilePin_355,profilePin_356,profilePin_357,profilePin_358,profilePin_359};
  wire  profilePin_360 = core__GEN_238_0;
  wire  profilePin_361 = core__GEN_239;
  wire  profilePin_362 = core__GEN_240_0;
  wire  profilePin_363 = core__GEN_241_0;
  wire  profilePin_364 = core__GEN_242;
  wire  profilePin_365 = core__GEN_243_0;
  wire  profilePin_366 = core__GEN_244_0;
  wire  profilePin_367 = core__GEN_245;
  wire  profilePin_368 = core__GEN_246_0;
  wire [369:0] _GEN_987 = {_GEN_978,profilePin_360,profilePin_361,profilePin_362,profilePin_363,profilePin_364,profilePin_365,profilePin_366,profilePin_367,profilePin_368};
  wire  profilePin_369 = core__GEN_247_0;
  wire  profilePin_370 = core__GEN_248_0;
  wire  profilePin_371 = core__GEN_249_0;
  wire  profilePin_372 = core__GEN_250_0;
  wire  profilePin_373 = core__GEN_251;
  wire  profilePin_374 = core__GEN_252_0;
  wire  profilePin_375 = core__GEN_253_0;
  wire  profilePin_376 = core__GEN_254;
  wire  profilePin_377 = core__GEN_255_0;
  wire [378:0] _GEN_996 = {_GEN_987,profilePin_369,profilePin_370,profilePin_371,profilePin_372,profilePin_373,profilePin_374,profilePin_375,profilePin_376,profilePin_377};
  wire  profilePin_378 = core__GEN_256_0;
  wire  profilePin_379 = core__GEN_257;
  wire  profilePin_380 = core__GEN_258_0;
  wire  profilePin_381 = core__GEN_259_0;
  wire  profilePin_382 = core__GEN_260;
  wire  profilePin_383 = core__GEN_261_0;
  wire  profilePin_384 = core__GEN_262_0;
  wire  profilePin_385 = core__GEN_263;
  wire  profilePin_386 = core__GEN_264_0;
  wire [387:0] _GEN_1005 = {_GEN_996,profilePin_378,profilePin_379,profilePin_380,profilePin_381,profilePin_382,profilePin_383,profilePin_384,profilePin_385,profilePin_386};
  wire  profilePin_387 = core__GEN_265_0;
  wire  profilePin_388 = core__GEN_266;
  wire  profilePin_389 = core__GEN_267_0;
  wire  profilePin_390 = core__GEN_268_0;
  wire  profilePin_391 = core__GEN_269;
  wire  profilePin_392 = core__GEN_270_0;
  wire  profilePin_393 = core__GEN_271_0;
  wire  profilePin_394 = core__GEN_272;
  wire  profilePin_395 = core__GEN_273_0;
  wire [396:0] _GEN_1014 = {_GEN_1005,profilePin_387,profilePin_388,profilePin_389,profilePin_390,profilePin_391,profilePin_392,profilePin_393,profilePin_394,profilePin_395};
  wire  profilePin_396 = core__GEN_274_0;
  wire  profilePin_397 = core__GEN_275;
  wire  profilePin_398 = core__GEN_276_0;
  wire  profilePin_399 = core__GEN_277_0;
  wire  profilePin_400 = core__GEN_278;
  wire  profilePin_401 = core__GEN_279;
  wire  profilePin_402 = core__GEN_280_0;
  wire  profilePin_403 = core__GEN_281;
  wire  profilePin_404 = core__GEN_282;
  wire [405:0] _GEN_1023 = {_GEN_1014,profilePin_396,profilePin_397,profilePin_398,profilePin_399,profilePin_400,profilePin_401,profilePin_402,profilePin_403,profilePin_404};
  wire  profilePin_405 = core__GEN_283_0;
  wire  profilePin_406 = core__GEN_284;
  wire  profilePin_407 = core__GEN_285;
  wire  profilePin_408 = core__GEN_286_0;
  wire  profilePin_409 = core__GEN_287;
  wire  profilePin_410 = core__GEN_288;
  wire  profilePin_411 = core__GEN_289_0;
  wire  profilePin_412 = core__GEN_290;
  wire  profilePin_413 = core__GEN_291;
  wire [414:0] _GEN_1032 = {_GEN_1023,profilePin_405,profilePin_406,profilePin_407,profilePin_408,profilePin_409,profilePin_410,profilePin_411,profilePin_412,profilePin_413};
  wire  profilePin_414 = core__GEN_292_0;
  wire  profilePin_415 = core__GEN_293_0;
  wire  profilePin_416 = core__GEN_294;
  wire  profilePin_417 = core__GEN_295_0;
  wire  profilePin_418 = core__GEN_296_0;
  wire  profilePin_419 = core__GEN_297_0;
  wire  profilePin_420 = core__GEN_298_0;
  wire  profilePin_421 = core__GEN_299_0;
  wire  profilePin_422 = core__GEN_300;
  wire [423:0] _GEN_1041 = {_GEN_1032,profilePin_414,profilePin_415,profilePin_416,profilePin_417,profilePin_418,profilePin_419,profilePin_420,profilePin_421,profilePin_422};
  wire  profilePin_423 = core__GEN_301_0;
  wire  profilePin_424 = core__GEN_302_0;
  wire  profilePin_425 = core__GEN_303_0;
  wire  profilePin_426 = core__GEN_304_0;
  wire  profilePin_427 = core__GEN_305_0;
  wire  profilePin_428 = core__GEN_306;
  wire  profilePin_429 = core__GEN_307_0;
  wire  profilePin_430 = core__GEN_308_0;
  wire  profilePin_431 = core__GEN_309_0;
  wire [432:0] _GEN_1050 = {_GEN_1041,profilePin_423,profilePin_424,profilePin_425,profilePin_426,profilePin_427,profilePin_428,profilePin_429,profilePin_430,profilePin_431};
  wire  profilePin_432 = core__GEN_310_0;
  wire  profilePin_433 = core__GEN_311_0;
  wire  profilePin_434 = core__GEN_312;
  wire  profilePin_435 = core__GEN_313_0;
  wire  profilePin_436 = core__GEN_314_0;
  wire  profilePin_437 = core__GEN_315_0;
  wire  profilePin_438 = core__GEN_316_0;
  wire  profilePin_439 = core__GEN_317;
  wire  profilePin_440 = core__GEN_318;
  wire [441:0] _GEN_1059 = {_GEN_1050,profilePin_432,profilePin_433,profilePin_434,profilePin_435,profilePin_436,profilePin_437,profilePin_438,profilePin_439,profilePin_440};
  wire  profilePin_441 = core__GEN_319_0;
  wire  profilePin_442 = core__GEN_320_0;
  wire  profilePin_443 = core__GEN_321_0;
  wire  profilePin_444 = core__GEN_322_0;
  wire  profilePin_445 = core__GEN_323;
  wire  profilePin_446 = core__GEN_324;
  wire  profilePin_447 = core__GEN_325;
  wire  profilePin_448 = core__GEN_326;
  wire  profilePin_449 = core__GEN_327;
  wire [450:0] _GEN_1068 = {_GEN_1059,profilePin_441,profilePin_442,profilePin_443,profilePin_444,profilePin_445,profilePin_446,profilePin_447,profilePin_448,profilePin_449};
  wire  profilePin_450 = core__GEN_328;
  wire  profilePin_451 = core__GEN_329;
  wire  profilePin_452 = core__GEN_330;
  wire  profilePin_453 = core__GEN_331;
  wire  profilePin_454 = core__GEN_332;
  wire  profilePin_455 = core__GEN_333;
  wire  profilePin_456 = core__GEN_334;
  wire  profilePin_457 = core__GEN_335;
  wire  profilePin_458 = core__GEN_336;
  wire [459:0] _GEN_1077 = {_GEN_1068,profilePin_450,profilePin_451,profilePin_452,profilePin_453,profilePin_454,profilePin_455,profilePin_456,profilePin_457,profilePin_458};
  wire  profilePin_459 = core__GEN_337;
  wire  profilePin_460 = core__GEN_338;
  wire  profilePin_461 = core__GEN_339;
  wire  profilePin_462 = core__GEN_340;
  wire  profilePin_463 = core__GEN_341;
  wire  profilePin_464 = core__GEN_342;
  wire  profilePin_465 = core__GEN_343;
  wire  profilePin_466 = core__GEN_344;
  wire  profilePin_467 = core__GEN_345;
  wire [468:0] _GEN_1086 = {_GEN_1077,profilePin_459,profilePin_460,profilePin_461,profilePin_462,profilePin_463,profilePin_464,profilePin_465,profilePin_466,profilePin_467};
  wire  profilePin_468 = core__GEN_346;
  wire  profilePin_469 = core__GEN_347;
  wire  profilePin_470 = core__GEN_348;
  wire  profilePin_471 = core__GEN_349;
  wire  profilePin_472 = core__GEN_350;
  wire  profilePin_473 = core__GEN_351;
  wire  profilePin_474 = core__GEN_352;
  wire  profilePin_475 = core__GEN_353;
  wire  profilePin_476 = core__GEN_354;
  wire [477:0] _GEN_1095 = {_GEN_1086,profilePin_468,profilePin_469,profilePin_470,profilePin_471,profilePin_472,profilePin_473,profilePin_474,profilePin_475,profilePin_476};
  wire  profilePin_477 = core__GEN_355;
  wire  profilePin_478 = core__GEN_356;
  wire  profilePin_479 = core__GEN_357;
  wire  profilePin_480 = core__GEN_358;
  wire  profilePin_481 = core__GEN_359;
  wire  profilePin_482 = core__GEN_360;
  wire  profilePin_483 = core__GEN_361;
  wire  profilePin_484 = core__GEN_362;
  wire  profilePin_485 = core__GEN_363;
  wire [486:0] _GEN_1104 = {_GEN_1095,profilePin_477,profilePin_478,profilePin_479,profilePin_480,profilePin_481,profilePin_482,profilePin_483,profilePin_484,profilePin_485};
  wire  profilePin_486 = core__GEN_364;
  wire  profilePin_487 = core__GEN_365;
  wire  profilePin_488 = core__GEN_366;
  wire  profilePin_489 = core__GEN_367;
  wire  profilePin_490 = core__GEN_368;
  wire  profilePin_491 = core__GEN_369;
  wire  profilePin_492 = core__GEN_370;
  wire  profilePin_493 = core__GEN_371;
  wire  profilePin_494 = core__GEN_372;
  wire [495:0] _GEN_1113 = {_GEN_1104,profilePin_486,profilePin_487,profilePin_488,profilePin_489,profilePin_490,profilePin_491,profilePin_492,profilePin_493,profilePin_494};
  wire  profilePin_495 = core__GEN_373;
  wire  profilePin_496 = core__GEN_374;
  wire  profilePin_497 = core__GEN_375;
  wire  profilePin_498 = core__GEN_376;
  wire  profilePin_499 = core__GEN_377;
  wire  profilePin_500 = core__GEN_378;
  wire  profilePin_501 = core__GEN_379;
  wire  profilePin_502 = core__GEN_380;
  wire  profilePin_503 = core__GEN_381;
  wire [504:0] _GEN_1122 = {_GEN_1113,profilePin_495,profilePin_496,profilePin_497,profilePin_498,profilePin_499,profilePin_500,profilePin_501,profilePin_502,profilePin_503};
  wire  profilePin_504 = core__GEN_382;
  wire  profilePin_505 = core__GEN_383;
  wire  profilePin_506 = core__GEN_384;
  wire  profilePin_507 = core__GEN_385;
  wire  profilePin_508 = core__GEN_386;
  wire  profilePin_509 = core__GEN_387;
  wire  profilePin_510 = core__GEN_388;
  wire  profilePin_511 = core__GEN_389;
  wire  profilePin_512 = core__GEN_390;
  wire [513:0] _GEN_1131 = {_GEN_1122,profilePin_504,profilePin_505,profilePin_506,profilePin_507,profilePin_508,profilePin_509,profilePin_510,profilePin_511,profilePin_512};
  wire  profilePin_513 = core__GEN_391;
  wire  profilePin_514 = core__GEN_392;
  wire  profilePin_515 = core__GEN_393;
  wire  profilePin_516 = core__GEN_394;
  wire  profilePin_517 = core__GEN_395;
  wire  profilePin_518 = core__GEN_396;
  wire  profilePin_519 = core__GEN_397;
  wire  profilePin_520 = core__GEN_398;
  wire  profilePin_521 = core__GEN_399;
  wire [522:0] _GEN_1140 = {_GEN_1131,profilePin_513,profilePin_514,profilePin_515,profilePin_516,profilePin_517,profilePin_518,profilePin_519,profilePin_520,profilePin_521};
  wire  profilePin_522 = core__GEN_400;
  wire  profilePin_523 = core__GEN_401;
  wire  profilePin_524 = core__GEN_402;
  wire  profilePin_525 = core__GEN_403;
  wire  profilePin_526 = core__GEN_404;
  wire  profilePin_527 = core__GEN_405;
  wire  profilePin_528 = core__GEN_406;
  wire  profilePin_529 = core__GEN_407;
  wire  profilePin_530 = core__GEN_408;
  wire [531:0] _GEN_1149 = {_GEN_1140,profilePin_522,profilePin_523,profilePin_524,profilePin_525,profilePin_526,profilePin_527,profilePin_528,profilePin_529,profilePin_530};
  wire  profilePin_531 = core__GEN_409;
  wire  profilePin_532 = core__GEN_410;
  wire  profilePin_533 = core__GEN_411;
  wire  profilePin_534 = core__GEN_412;
  wire  profilePin_535 = core__GEN_413;
  wire  profilePin_536 = core__GEN_414;
  wire  profilePin_537 = core__GEN_415;
  wire  profilePin_538 = core__GEN_416;
  wire  profilePin_539 = core__GEN_417;
  wire [540:0] _GEN_1158 = {_GEN_1149,profilePin_531,profilePin_532,profilePin_533,profilePin_534,profilePin_535,profilePin_536,profilePin_537,profilePin_538,profilePin_539};
  wire  profilePin_540 = core__GEN_418;
  wire  profilePin_541 = core__GEN_419;
  wire  profilePin_542 = core__GEN_420;
  wire  profilePin_543 = core__GEN_421;
  wire  profilePin_544 = core__GEN_422;
  wire  profilePin_545 = core__GEN_423;
  wire  profilePin_546 = core__GEN_424;
  wire  profilePin_547 = core__GEN_425;
  wire  profilePin_548 = core__GEN_426;
  wire [549:0] _GEN_1167 = {_GEN_1158,profilePin_540,profilePin_541,profilePin_542,profilePin_543,profilePin_544,profilePin_545,profilePin_546,profilePin_547,profilePin_548};
  wire  profilePin_549 = core__GEN_427;
  wire  profilePin_550 = core__GEN_428;
  wire  profilePin_551 = core__GEN_429;
  wire  profilePin_552 = core__GEN_430;
  wire  profilePin_553 = core__GEN_431;
  wire  profilePin_554 = core__GEN_432;
  wire  profilePin_555 = core__GEN_433;
  wire  profilePin_556 = core__GEN_434;
  wire  profilePin_557 = core__GEN_435;
  wire [558:0] _GEN_1176 = {_GEN_1167,profilePin_549,profilePin_550,profilePin_551,profilePin_552,profilePin_553,profilePin_554,profilePin_555,profilePin_556,profilePin_557};
  wire  profilePin_558 = core__GEN_436;
  wire  profilePin_559 = core__GEN_437;
  wire  profilePin_560 = core__GEN_438;
  wire  profilePin_561 = core__GEN_439;
  wire  profilePin_562 = core__GEN_440;
  wire  profilePin_563 = core__GEN_441;
  wire  profilePin_564 = core__GEN_442;
  wire  profilePin_565 = core__GEN_443;
  wire  profilePin_566 = core__GEN_444;
  wire [567:0] _GEN_1185 = {_GEN_1176,profilePin_558,profilePin_559,profilePin_560,profilePin_561,profilePin_562,profilePin_563,profilePin_564,profilePin_565,profilePin_566};
  wire  profilePin_567 = core__GEN_445;
  wire  profilePin_568 = core__GEN_446;
  wire  profilePin_569 = core__GEN_447;
  wire  profilePin_570 = core__GEN_448;
  wire  profilePin_571 = core__GEN_449;
  wire  profilePin_572 = core__GEN_450;
  wire  profilePin_573 = core__GEN_451;
  wire  profilePin_574 = core__GEN_452;
  wire  profilePin_575 = core__GEN_453;
  wire [576:0] _GEN_1194 = {_GEN_1185,profilePin_567,profilePin_568,profilePin_569,profilePin_570,profilePin_571,profilePin_572,profilePin_573,profilePin_574,profilePin_575};
  wire  profilePin_576 = core__GEN_454;
  wire  profilePin_577 = core__GEN_455;
  wire  profilePin_578 = core__GEN_456;
  wire  profilePin_579 = core__GEN_457;
  wire  profilePin_580 = core__GEN_458;
  wire  profilePin_581 = core__GEN_459;
  wire  profilePin_582 = core__GEN_460;
  wire  profilePin_583 = core__GEN_461;
  wire  profilePin_584 = core__GEN_462;
  wire [585:0] _GEN_1203 = {_GEN_1194,profilePin_576,profilePin_577,profilePin_578,profilePin_579,profilePin_580,profilePin_581,profilePin_582,profilePin_583,profilePin_584};
  wire  profilePin_586 = core__GEN_0;
  wire  profilePin_587 = core__GEN_1_2;
  wire  profilePin_588 = core__GEN_2;
  wire  profilePin_589 = core__GEN_3;
  wire  profilePin_590 = core__GEN_4_1;
  wire  profilePin_591 = core__GEN_5;
  wire  profilePin_592 = core__GEN_6;
  wire  profilePin_593 = core__GEN_7_1;
  wire  profilePin_594 = core__GEN_8;
  wire [594:0] _GEN_1212 = {_GEN_1203,profilePin_586,profilePin_587,profilePin_588,profilePin_589,profilePin_590,profilePin_591,profilePin_592,profilePin_593,profilePin_594};
  wire  profilePin_595 = core__GEN_9;
  wire  profilePin_596 = core__GEN_10_2;
  wire  profilePin_597 = core__GEN_11;
  wire  profilePin_598 = core__GEN_12;
  wire  profilePin_599 = core__GEN_13_1;
  wire  profilePin_600 = core__GEN_14_0;
  wire  profilePin_601 = core__GEN_15_1;
  wire  profilePin_602 = core__GEN_16_0;
  wire  profilePin_603 = core__GEN_17_1;
  wire [603:0] _GEN_1221 = {_GEN_1212,profilePin_595,profilePin_596,profilePin_597,profilePin_598,profilePin_599,profilePin_600,profilePin_601,profilePin_602,profilePin_603};
  wire  profilePin_604 = core__GEN_18_1;
  wire  profilePin_605 = core__GEN_19;
  wire  profilePin_606 = core__GEN_20;
  wire  profilePin_607 = core__GEN_21;
  wire  profilePin_608 = core__GEN_22;
  wire  profilePin_609 = core__GEN_23;
  wire  profilePin_610 = memory__GEN_0_1;
  wire  profilePin_611 = memory__GEN_1_0;
  wire  profilePin_612 = memory__GEN_2_1;
  wire [612:0] _GEN_1230 = {_GEN_1221,profilePin_604,profilePin_605,profilePin_606,profilePin_607,profilePin_608,profilePin_609,profilePin_610,profilePin_611,profilePin_612};
  wire  profilePin_613 = memory__GEN_3_1;
  wire  profilePin_614 = memory__GEN_4_0;
  wire [614:0] _GEN_1232 = {_GEN_1230,profilePin_613,profilePin_614};
  wire  profilePin_615 = memory__GEN_5_1;
  Core core ( // @[top.scala 26:26]
    .metaReset(core_metaReset),
    .clock(core_clock),
    .reset(core_reset),
    .io_imem_req_bits_addr(core_io_imem_req_bits_addr),
    .io_imem_resp_bits_data(core_io_imem_resp_bits_data),
    .io_dmem_req_bits_addr(core_io_dmem_req_bits_addr),
    .io_dmem_req_bits_data(core_io_dmem_req_bits_data),
    .io_dmem_req_bits_fcn(core_io_dmem_req_bits_fcn),
    .io_dmem_req_bits_typ(core_io_dmem_req_bits_typ),
    .io_dmem_resp_bits_data(core_io_dmem_resp_bits_data),
    ._GEN_411(core__GEN_411),
    ._GEN_405(core__GEN_405),
    ._GEN_92(core__GEN_92),
    ._GEN_52(core__GEN_52),
    ._GEN_305(core__GEN_305),
    ._GEN_200(core__GEN_200),
    ._GEN_149(core__GEN_149),
    ._GEN_426(core__GEN_426),
    ._GEN_291(core__GEN_291),
    ._GEN_1_0(core__GEN_1_0),
    ._GEN_25(core__GEN_25),
    ._GEN_248(core__GEN_248),
    ._GEN_107(core__GEN_107),
    ._GEN_134(core__GEN_134),
    ._GEN_206(core__GEN_206),
    ._GEN_40(core__GEN_40),
    ._GEN_306(core__GEN_306),
    ._GEN_233(core__GEN_233),
    ._GEN_128(core__GEN_128),
    ._GEN_384(core__GEN_384),
    ._GEN_191(core__GEN_191),
    ._GEN_16(core__GEN_16),
    ._GEN_227(core__GEN_227),
    ._GEN_19(core__GEN_19),
    ._GEN_327(core__GEN_327),
    ._GEN_113(core__GEN_113),
    ._GEN_46(core__GEN_46),
    ._GEN_299(core__GEN_299),
    ._GEN_390(core__GEN_390),
    ._GEN_73(core__GEN_73),
    ._GEN_212(core__GEN_212),
    ._GEN_10(core__GEN_10),
    ._GEN_285(core__GEN_285),
    ._GEN_318(core__GEN_318),
    ._GEN_312(core__GEN_312),
    ._GEN_31(core__GEN_31),
    ._GEN_311(core__GEN_311),
    ._GEN_67(core__GEN_67),
    ._GEN_320(core__GEN_320),
    ._GEN_399(core__GEN_399),
    ._GEN_215(core__GEN_215),
    ._GEN_221(core__GEN_221),
    ._GEN_101(core__GEN_101),
    ._GEN_110(core__GEN_110),
    ._GEN_387(core__GEN_387),
    ._GEN_283(core__GEN_283),
    ._GEN_314(core__GEN_314),
    ._GEN_178(core__GEN_178),
    ._GEN_209(core__GEN_209),
    ._GEN_300(core__GEN_300),
    ._GEN_279(core__GEN_279),
    ._GEN_269(core__GEN_269),
    ._GEN_28(core__GEN_28),
    ._GEN_277(core__GEN_277),
    ._GEN_378(core__GEN_378),
    ._GEN_368(core__GEN_368),
    ._GEN_55(core__GEN_55),
    ._GEN_377(core__GEN_377),
    ._GEN_194(core__GEN_194),
    ._GEN_22(core__GEN_22),
    ._GEN_12(core__GEN_12),
    ._GEN_294(core__GEN_294),
    ._GEN_13(core__GEN_13),
    ._GEN_49(core__GEN_49),
    ._GEN_116(core__GEN_116),
    ._GEN_393(core__GEN_393),
    ._GEN_362(core__GEN_362),
    ._GEN_7(core__GEN_7),
    ._GEN_461(core__GEN_461),
    ._GEN_34(core__GEN_34),
    ._GEN_122(core__GEN_122),
    ._GEN_308(core__GEN_308),
    ._GEN_263(core__GEN_263),
    ._GEN_95(core__GEN_95),
    ._GEN_230(core__GEN_230),
    ._GEN_293(core__GEN_293),
    ._GEN_184(core__GEN_184),
    ._GEN_1_1(core__GEN_1_1),
    ._GEN_10_0(core__GEN_10_0),
    ._GEN_197(core__GEN_197),
    ._GEN_187(core__GEN_187),
    ._GEN_449(core__GEN_449),
    ._GEN_288(core__GEN_288),
    ._GEN_104(core__GEN_104),
    ._GEN_265(core__GEN_265),
    ._GEN_296(core__GEN_296),
    ._GEN_160(core__GEN_160),
    ._GEN_172(core__GEN_172),
    ._GEN_203(core__GEN_203),
    ._GEN_245(core__GEN_245),
    ._GEN_0(core__GEN_0),
    ._GEN_272(core__GEN_272),
    ._GEN_271(core__GEN_271),
    ._GEN_37(core__GEN_37),
    ._GEN_166(core__GEN_166),
    ._GEN_280(core__GEN_280),
    ._GEN_286(core__GEN_286),
    ._GEN_381(core__GEN_381),
    ._GEN_371(core__GEN_371),
    ._GEN_266(core__GEN_266),
    ._GEN_16_0(core__GEN_16_0),
    ._GEN_22_0(core__GEN_22_0),
    ._GEN_302(core__GEN_302),
    ._GEN_344(core__GEN_344),
    ._GEN_282(core__GEN_282),
    ._GEN_443(core__GEN_443),
    ._GEN_16_1(core__GEN_16_1),
    ._GEN_251(core__GEN_251),
    ._GEN_10_1(core__GEN_10_1),
    ._GEN_259(core__GEN_259),
    ._GEN_98(core__GEN_98),
    ._GEN_6(core__GEN_6),
    ._GEN_350(core__GEN_350),
    ._GEN_365(core__GEN_365),
    ._GEN_15(core__GEN_15),
    ._GEN_152(core__GEN_152),
    ._GEN_446(core__GEN_446),
    ._GEN_332(core__GEN_332),
    ._GEN_326(core__GEN_326),
    ._GEN_19_0(core__GEN_19_0),
    ._GEN_148(core__GEN_148),
    ._GEN_359(core__GEN_359),
    ._GEN_15_0(core__GEN_15_0),
    ._GEN_87(core__GEN_87),
    ._GEN_458(core__GEN_458),
    ._GEN_452(core__GEN_452),
    ._GEN_13_0(core__GEN_13_0),
    ._GEN_3(core__GEN_3),
    ._GEN_347(core__GEN_347),
    ._GEN_274(core__GEN_274),
    ._GEN_425(core__GEN_425),
    ._GEN_239(core__GEN_239),
    ._GEN_232(core__GEN_232),
    ._GEN_190(core__GEN_190),
    ._GEN_154(core__GEN_154),
    ._GEN_289(core__GEN_289),
    ._GEN_431(core__GEN_431),
    ._GEN_181(core__GEN_181),
    ._GEN_253(core__GEN_253),
    ._GEN_254(core__GEN_254),
    ._GEN_353(core__GEN_353),
    ._GEN_72(core__GEN_72),
    ._GEN_175(core__GEN_175),
    ._GEN_169(core__GEN_169),
    ._GEN_260(core__GEN_260),
    ._GEN_4_0(core__GEN_4_0),
    ._GEN_275(core__GEN_275),
    ._GEN_247(core__GEN_247),
    ._GEN_268(core__GEN_268),
    ._GEN_9(core__GEN_9),
    ._GEN_338(core__GEN_338),
    ._GEN_374(core__GEN_374),
    ._GEN_242(core__GEN_242),
    ._GEN_214(core__GEN_214),
    ._GEN_250(core__GEN_250),
    ._GEN_455(core__GEN_455),
    ._GEN_241(core__GEN_241),
    ._GEN_142(core__GEN_142),
    ._GEN_136(core__GEN_136),
    ._GEN_413(core__GEN_413),
    ._GEN_235(core__GEN_235),
    ._GEN_236(core__GEN_236),
    ._GEN_262(core__GEN_262),
    ._GEN_335(core__GEN_335),
    ._GEN_54(core__GEN_54),
    ._GEN_313(core__GEN_313),
    ._GEN_18(core__GEN_18),
    ._GEN_69(core__GEN_69),
    ._GEN_157(core__GEN_157),
    ._GEN_434(core__GEN_434),
    ._GEN_248_0(core__GEN_248_0),
    ._GEN_257(core__GEN_257),
    ._GEN_320_0(core__GEN_320_0),
    ._GEN_75(core__GEN_75),
    ._GEN_356(core__GEN_356),
    ._GEN_12_0(core__GEN_12_0),
    ._GEN_90(core__GEN_90),
    ._GEN_163(core__GEN_163),
    ._GEN_419(core__GEN_419),
    ._GEN_314_0(core__GEN_314_0),
    ._GEN_7_0(core__GEN_7_0),
    ._GEN_130(core__GEN_130),
    ._GEN_341(core__GEN_341),
    ._GEN_440(core__GEN_440),
    ._GEN_229(core__GEN_229),
    ._GEN_299_0(core__GEN_299_0),
    ._GEN_121(core__GEN_121),
    ._GEN_256(core__GEN_256),
    ._GEN_398(core__GEN_398),
    ._GEN_81(core__GEN_81),
    ._GEN_407(core__GEN_407),
    ._GEN_149_0(core__GEN_149_0),
    ._GEN_416(core__GEN_416),
    ._GEN_281(core__GEN_281),
    ._GEN_15_1(core__GEN_15_1),
    ._GEN_380(core__GEN_380),
    ._GEN_57(core__GEN_57),
    ._GEN_145(core__GEN_145),
    ._GEN_296_0(core__GEN_296_0),
    ._GEN_223(core__GEN_223),
    ._GEN_118(core__GEN_118),
    ._GEN_322(core__GEN_322),
    ._GEN_422(core__GEN_422),
    ._GEN_244(core__GEN_244),
    ._GEN_124(core__GEN_124),
    ._GEN_103(core__GEN_103),
    ._GEN_238(core__GEN_238),
    ._GEN_329(core__GEN_329),
    ._GEN_63(core__GEN_63),
    ._GEN_151(core__GEN_151),
    ._GEN_202(core__GEN_202),
    ._GEN_6_0(core__GEN_6_0),
    ._GEN_196(core__GEN_196),
    ._GEN_437(core__GEN_437),
    ._GEN_302_0(core__GEN_302_0),
    ._GEN_295(core__GEN_295),
    ._GEN_301(core__GEN_301),
    ._GEN_310(core__GEN_310),
    ._GEN_401(core__GEN_401),
    ._GEN_395(core__GEN_395),
    ._GEN_78(core__GEN_78),
    ._GEN_84(core__GEN_84),
    ._GEN_217(core__GEN_217),
    ._GEN_428(core__GEN_428),
    ._GEN_308_0(core__GEN_308_0),
    ._GEN_323(core__GEN_323),
    ._GEN_36(core__GEN_36),
    ._GEN_42(core__GEN_42),
    ._GEN_317(core__GEN_317),
    ._GEN_316(core__GEN_316),
    ._GEN_139(core__GEN_139),
    ._GEN_404(core__GEN_404),
    ._GEN_290(core__GEN_290),
    ._GEN_18_0(core__GEN_18_0),
    ._GEN_226(core__GEN_226),
    ._GEN_106(core__GEN_106),
    ._GEN_51(core__GEN_51),
    ._GEN_45(core__GEN_45),
    ._GEN_9_0(core__GEN_9_0),
    ._GEN_367(core__GEN_367),
    ._GEN_319(core__GEN_319),
    ._GEN_284(core__GEN_284),
    ._GEN_274_0(core__GEN_274_0),
    ._GEN_39(core__GEN_39),
    ._GEN_383(core__GEN_383),
    ._GEN_373(core__GEN_373),
    ._GEN_66(core__GEN_66),
    ._GEN_18_1(core__GEN_18_1),
    ._GEN_410(core__GEN_410),
    ._GEN_24(core__GEN_24),
    ._GEN_305_0(core__GEN_305_0),
    ._GEN_112(core__GEN_112),
    ._GEN_211(core__GEN_211),
    ._GEN_220(core__GEN_220),
    ._GEN_8(core__GEN_8),
    ._GEN_2(core__GEN_2),
    ._GEN_311_0(core__GEN_311_0),
    ._GEN_133(core__GEN_133),
    ._GEN_127(core__GEN_127),
    ._GEN_288_0(core__GEN_288_0),
    ._GEN_389(core__GEN_389),
    ._GEN_91(core__GEN_91),
    ._GEN_205(core__GEN_205),
    ._GEN_100(core__GEN_100),
    ._GEN_304(core__GEN_304),
    ._GEN_60(core__GEN_60),
    ._GEN_298(core__GEN_298),
    ._GEN_189(core__GEN_189),
    ._GEN_199(core__GEN_199),
    ._GEN_177(core__GEN_177),
    ._GEN_12_1(core__GEN_12_1),
    ._GEN_268_0(core__GEN_268_0),
    ._GEN_94(core__GEN_94),
    ._GEN_376(core__GEN_376),
    ._GEN_162(core__GEN_162),
    ._GEN_193(core__GEN_193),
    ._GEN_208(core__GEN_208),
    ._GEN_454(core__GEN_454),
    ._GEN_293_0(core__GEN_293_0),
    ._GEN_261(core__GEN_261),
    ._GEN_115(core__GEN_115),
    ._GEN_27(core__GEN_27),
    ._GEN_270(core__GEN_270),
    ._GEN_392(core__GEN_392),
    ._GEN_361(core__GEN_361),
    ._GEN_287(core__GEN_287),
    ._GEN_183(core__GEN_183),
    ._GEN_256_0(core__GEN_256_0),
    ._GEN_460(core__GEN_460),
    ._GEN_278(core__GEN_278),
    ._GEN_33(core__GEN_33),
    ._GEN_276(core__GEN_276),
    ._GEN_282_0(core__GEN_282_0),
    ._GEN_292(core__GEN_292),
    ._GEN_355(core__GEN_355),
    ._GEN_48(core__GEN_48),
    ._GEN_386(core__GEN_386),
    ._GEN_6_1(core__GEN_6_1),
    ._GEN_277_0(core__GEN_277_0),
    ._GEN_21(core__GEN_21),
    ._GEN_307(core__GEN_307),
    ._GEN_262_0(core__GEN_262_0),
    ._GEN_109(core__GEN_109),
    ._GEN_11(core__GEN_11),
    ._GEN_244_0(core__GEN_244_0),
    ._GEN_448(core__GEN_448),
    ._GEN_442(core__GEN_442),
    ._GEN_21_0(core__GEN_21_0),
    ._GEN_15_2(core__GEN_15_2),
    ._GEN_457(core__GEN_457),
    ._GEN_337(core__GEN_337),
    ._GEN_30(core__GEN_30),
    ._GEN_83(core__GEN_83),
    ._GEN_364(core__GEN_364),
    ._GEN_171(core__GEN_171),
    ._GEN_186(core__GEN_186),
    ._GEN_328(core__GEN_328),
    ._GEN_463(core__GEN_463),
    ._GEN_144(core__GEN_144),
    ._GEN_279_0(core__GEN_279_0),
    ._GEN_436(core__GEN_436),
    ._GEN_97(core__GEN_97),
    ._GEN_9_1(core__GEN_9_1),
    ._GEN_264(core__GEN_264),
    ._GEN_165(core__GEN_165),
    ._GEN_159(core__GEN_159),
    ._GEN_370(core__GEN_370),
    ._GEN_250_0(core__GEN_250_0),
    ._GEN_265_0(core__GEN_265_0),
    ._GEN_258(core__GEN_258),
    ._GEN_5(core__GEN_5),
    ._GEN_285_0(core__GEN_285_0),
    ._GEN_180(core__GEN_180),
    ._GEN_271_0(core__GEN_271_0),
    ._GEN_9_2(core__GEN_9_2),
    ._GEN_243(core__GEN_243),
    ._GEN_349(core__GEN_349),
    ._GEN_343(core__GEN_343),
    ._GEN_147(core__GEN_147),
    ._GEN_77(core__GEN_77),
    ._GEN_352(core__GEN_352),
    ._GEN_174(core__GEN_174),
    ._GEN_225(core__GEN_225),
    ._GEN_247_0(core__GEN_247_0),
    ._GEN_252(core__GEN_252),
    ._GEN_325(core__GEN_325),
    ._GEN_132(core__GEN_132),
    ._GEN_147_0(core__GEN_147_0),
    ._GEN_151_0(core__GEN_151_0),
    ._GEN_238_0(core__GEN_238_0),
    ._GEN_240(core__GEN_240),
    ._GEN_451(core__GEN_451),
    ._GEN_65(core__GEN_65),
    ._GEN_273(core__GEN_273),
    ._GEN_346(core__GEN_346),
    ._GEN_59(core__GEN_59),
    ._GEN_409(core__GEN_409),
    ._GEN_231(core__GEN_231),
    ._GEN_253_0(core__GEN_253_0),
    ._GEN_331(core__GEN_331),
    ._GEN_86(core__GEN_86),
    ._GEN_8_0(core__GEN_8_0),
    ._GEN_80(core__GEN_80),
    ._GEN_11_0(core__GEN_11_0),
    ._GEN_430(core__GEN_430),
    ._GEN_424(core__GEN_424),
    ._GEN_3_1(core__GEN_3_1),
    ._GEN_246(core__GEN_246),
    ._GEN_12_2(core__GEN_12_2),
    ._GEN_71(core__GEN_71),
    ._GEN_153(core__GEN_153),
    ._GEN_168(core__GEN_168),
    ._GEN_445(core__GEN_445),
    ._GEN_310_0(core__GEN_310_0),
    ._GEN_259_0(core__GEN_259_0),
    ._GEN_267(core__GEN_267),
    ._GEN_126(core__GEN_126),
    ._GEN_358(core__GEN_358),
    ._GEN_213(core__GEN_213),
    ._GEN_255(core__GEN_255),
    ._GEN_334(core__GEN_334),
    ._GEN_156(core__GEN_156),
    ._GEN_150(core__GEN_150),
    ._GEN_412(core__GEN_412),
    ._GEN_114(core__GEN_114),
    ._GEN_228(core__GEN_228),
    ._GEN_141(core__GEN_141),
    ._GEN_11_1(core__GEN_11_1),
    ._GEN_418(core__GEN_418),
    ._GEN_427(core__GEN_427),
    ._GEN_313_0(core__GEN_313_0),
    ._GEN_292_0(core__GEN_292_0),
    ._GEN_241_0(core__GEN_241_0),
    ._GEN_108(core__GEN_108),
    ._GEN_249(core__GEN_249),
    ._GEN_6_2(core__GEN_6_2),
    ._GEN_340(core__GEN_340),
    ._GEN_312_0(core__GEN_312_0),
    ._GEN_68(core__GEN_68),
    ._GEN_74(core__GEN_74),
    ._GEN_207(core__GEN_207),
    ._GEN_235_0(core__GEN_235_0),
    ._GEN_439(core__GEN_439),
    ._GEN_20(core__GEN_20),
    ._GEN_298_0(core__GEN_298_0),
    ._GEN_307_0(core__GEN_307_0),
    ._GEN_234(core__GEN_234),
    ._GEN_306_0(core__GEN_306_0),
    ._GEN_129(core__GEN_129),
    ._GEN_17(core__GEN_17),
    ._GEN_406(core__GEN_406),
    ._GEN_89(core__GEN_89),
    ._GEN_433(core__GEN_433),
    ._GEN_319_0(core__GEN_319_0),
    ._GEN_47(core__GEN_47),
    ._GEN_53(core__GEN_53),
    ._GEN_135(core__GEN_135),
    ._GEN_391(core__GEN_391),
    ._GEN_400(core__GEN_400),
    ._GEN_415(core__GEN_415),
    ._GEN_222(core__GEN_222),
    ._GEN_295_0(core__GEN_295_0),
    ._GEN_270_0(core__GEN_270_0),
    ._GEN_29(core__GEN_29),
    ._GEN_4_1(core__GEN_4_1),
    ._GEN_322_0(core__GEN_322_0),
    ._GEN_41(core__GEN_41),
    ._GEN_56(core__GEN_56),
    ._GEN_14(core__GEN_14),
    ._GEN_195(core__GEN_195),
    ._GEN_421(core__GEN_421),
    ._GEN_280_0(core__GEN_280_0),
    ._GEN_237(core__GEN_237),
    ._GEN_102(core__GEN_102),
    ._GEN_379(core__GEN_379),
    ._GEN_62(core__GEN_62),
    ._GEN_394(core__GEN_394),
    ._GEN_23(core__GEN_23),
    ._GEN_35(core__GEN_35),
    ._GEN_123(core__GEN_123),
    ._GEN_117(core__GEN_117),
    ._GEN_369(core__GEN_369),
    ._GEN_321(core__GEN_321),
    ._GEN_216(core__GEN_216),
    ._GEN_5_1(core__GEN_5_1),
    ._GEN_14_0(core__GEN_14_0),
    ._GEN_13_1(core__GEN_13_1),
    ._GEN_316_0(core__GEN_316_0),
    ._GEN_294_0(core__GEN_294_0),
    ._GEN_50(core__GEN_50),
    ._GEN_138(core__GEN_138),
    ._GEN_201(core__GEN_201),
    ._GEN_210(core__GEN_210),
    ._GEN_96(core__GEN_96),
    ._GEN_301_0(core__GEN_301_0),
    ._GEN_315(core__GEN_315),
    ._GEN_309(core__GEN_309),
    ._GEN_17_0(core__GEN_17_0),
    ._GEN_283_0(core__GEN_283_0),
    ._GEN_273_0(core__GEN_273_0),
    ._GEN_105(core__GEN_105),
    ._GEN_382(core__GEN_382),
    ._GEN_303(core__GEN_303),
    ._GEN_204(core__GEN_204),
    ._GEN_318_0(core__GEN_318_0),
    ._GEN_173(core__GEN_173),
    ._GEN_198(core__GEN_198),
    ._GEN_258_0(core__GEN_258_0),
    ._GEN_304_0(core__GEN_304_0),
    ._GEN_23_0(core__GEN_23_0),
    ._GEN_272_0(core__GEN_272_0),
    ._GEN_120(core__GEN_120),
    ._GEN_403(core__GEN_403),
    ._GEN_372(core__GEN_372),
    ._GEN_366(core__GEN_366),
    ._GEN_267_0(core__GEN_267_0),
    ._GEN_188(core__GEN_188),
    ._GEN_289_0(core__GEN_289_0),
    ._GEN_1_2(core__GEN_1_2),
    ._GEN_44(core__GEN_44),
    ._GEN_287_0(core__GEN_287_0),
    ._GEN_297(core__GEN_297),
    ._GEN_388(core__GEN_388),
    ._GEN_397(core__GEN_397),
    ._GEN_2_1(core__GEN_2_1),
    ._GEN_252_0(core__GEN_252_0),
    ._GEN_450(core__GEN_450),
    ._GEN_99(core__GEN_99),
    ._GEN_351(core__GEN_351),
    ._GEN_38(core__GEN_38),
    ._GEN_111(core__GEN_111),
    ._GEN_219(core__GEN_219),
    ._GEN_17_1(core__GEN_17_1),
    ._GEN_7_1(core__GEN_7_1),
    ._GEN_453(core__GEN_453),
    ._GEN_447(core__GEN_447),
    ._GEN_26(core__GEN_26),
    ._GEN_176(core__GEN_176),
    ._GEN_182(core__GEN_182),
    ._GEN_438(core__GEN_438),
    ._GEN_333(core__GEN_333),
    ._GEN_290_0(core__GEN_290_0),
    ._GEN_240_0(core__GEN_240_0),
    ._GEN_0_1(core__GEN_0_1),
    ._GEN_339(core__GEN_339),
    ._GEN_32(core__GEN_32),
    ._GEN_161(core__GEN_161),
    ._GEN_275_0(core__GEN_275_0),
    ._GEN_170(core__GEN_170),
    ._GEN_375(core__GEN_375),
    ._GEN_261_0(core__GEN_261_0),
    ._GEN_192(core__GEN_192),
    ._GEN_20_0(core__GEN_20_0),
    ._GEN_255_0(core__GEN_255_0),
    ._GEN_269_0(core__GEN_269_0),
    ._GEN_10_2(core__GEN_10_2),
    ._GEN_360(core__GEN_360),
    ._GEN_281_0(core__GEN_281_0),
    ._GEN_291_0(core__GEN_291_0),
    ._GEN_155(core__GEN_155),
    ._GEN_88(core__GEN_88),
    ._GEN_300_0(core__GEN_300_0),
    ._GEN_432(core__GEN_432),
    ._GEN_11_2(core__GEN_11_2),
    ._GEN_286_0(core__GEN_286_0),
    ._GEN_276_0(core__GEN_276_0),
    ._GEN_5_2(core__GEN_5_2),
    ._GEN_254_0(core__GEN_254_0),
    ._GEN_93(core__GEN_93),
    ._GEN_5_3(core__GEN_5_3),
    ._GEN_459(core__GEN_459),
    ._GEN_385(core__GEN_385),
    ._GEN_354(core__GEN_354),
    ._GEN_234_0(core__GEN_234_0),
    ._GEN_3_2(core__GEN_3_2),
    ._GEN_146(core__GEN_146),
    ._GEN_441(core__GEN_441),
    ._GEN_321_0(core__GEN_321_0),
    ._GEN_14_1(core__GEN_14_1),
    ._GEN_257_0(core__GEN_257_0),
    ._GEN_13_2(core__GEN_13_2),
    ._GEN_348(core__GEN_348),
    ._GEN_82(core__GEN_82),
    ._GEN_357(core__GEN_357),
    ._GEN_243_0(core__GEN_243_0),
    ._GEN_8_1(core__GEN_8_1),
    ._GEN_8_2(core__GEN_8_2),
    ._GEN_462(core__GEN_462),
    ._GEN_456(core__GEN_456),
    ._GEN_342(core__GEN_342),
    ._GEN_278_0(core__GEN_278_0),
    ._GEN_70(core__GEN_70),
    ._GEN_158(core__GEN_158),
    ._GEN_420(core__GEN_420),
    ._GEN_414(core__GEN_414),
    ._GEN_236_0(core__GEN_236_0),
    ._GEN_185(core__GEN_185),
    ._GEN_336(core__GEN_336),
    ._GEN_61(core__GEN_61),
    ._GEN_143(core__GEN_143),
    ._GEN_284_0(core__GEN_284_0),
    ._GEN_179(core__GEN_179),
    ._GEN_435(core__GEN_435),
    ._GEN_242_0(core__GEN_242_0),
    ._GEN_249_0(core__GEN_249_0),
    ._GEN_137(core__GEN_137),
    ._GEN_76(core__GEN_76),
    ._GEN_164(core__GEN_164),
    ._GEN_237_0(core__GEN_237_0),
    ._GEN_315_0(core__GEN_315_0),
    ._GEN_264_0(core__GEN_264_0),
    ._GEN_263_0(core__GEN_263_0),
    ._GEN_363(core__GEN_363),
    ._GEN_167(core__GEN_167),
    ._GEN_246_0(core__GEN_246_0),
    ._GEN_43(core__GEN_43),
    ._GEN_266_0(core__GEN_266_0),
    ._GEN_131(core__GEN_131),
    ._GEN_125(core__GEN_125),
    ._GEN_317_0(core__GEN_317_0),
    ._GEN_224(core__GEN_224),
    ._GEN_150_0(core__GEN_150_0),
    ._GEN_119(core__GEN_119),
    ._GEN_239_0(core__GEN_239_0),
    ._GEN_330(core__GEN_330),
    ._GEN_152_0(core__GEN_152_0),
    ._GEN_146_0(core__GEN_146_0),
    ._GEN_7_2(core__GEN_7_2),
    ._GEN_297_0(core__GEN_297_0),
    ._GEN_245_0(core__GEN_245_0),
    ._GEN_11_3(core__GEN_11_3),
    ._GEN_345(core__GEN_345),
    ._GEN_323_0(core__GEN_323_0),
    ._GEN_396(core__GEN_396),
    ._GEN_79(core__GEN_79),
    ._GEN_218(core__GEN_218),
    ._GEN_408(core__GEN_408),
    ._GEN_423(core__GEN_423),
    ._GEN_309_0(core__GEN_309_0),
    ._GEN_303_0(core__GEN_303_0),
    ._GEN_64(core__GEN_64),
    ._GEN_417(core__GEN_417),
    ._GEN_429(core__GEN_429),
    ._GEN_444(core__GEN_444),
    ._GEN_324(core__GEN_324),
    ._GEN_58(core__GEN_58),
    ._GEN_251_0(core__GEN_251_0),
    ._GEN_260_0(core__GEN_260_0),
    ._GEN_140(core__GEN_140),
    ._GEN_402(core__GEN_402),
    ._GEN_85(core__GEN_85)
  );
  SyncScratchPadMemory memory ( // @[top.scala 29:28]
    .metaReset(memory_metaReset),
    .clock(memory_clock),
    .io_core_ports_0_req_bits_addr(memory_io_core_ports_0_req_bits_addr),
    .io_core_ports_0_req_bits_data(memory_io_core_ports_0_req_bits_data),
    .io_core_ports_0_req_bits_fcn(memory_io_core_ports_0_req_bits_fcn),
    .io_core_ports_0_req_bits_typ(memory_io_core_ports_0_req_bits_typ),
    .io_core_ports_0_resp_bits_data(memory_io_core_ports_0_resp_bits_data),
    ._GEN_1_0(memory__GEN_1_0),
    ._GEN_4_0(memory__GEN_4_0),
    ._GEN_0_1(memory__GEN_0_1),
    ._GEN_3_1(memory__GEN_3_1),
    ._GEN_2_1(memory__GEN_2_1),
    ._GEN_5_1(memory__GEN_5_1)
  );
  assign core_metaReset = metaReset;
  assign memory_metaReset = metaReset;
  assign io_imem_req_valid = 1'h1; // @[top.scala 34:22]
  assign io_imem_req_bits_addr = core_io_imem_req_bits_addr; // @[top.scala 34:22]
  assign io_imem_req_bits_data = 32'h0; // @[top.scala 34:22]
  assign io_imem_req_bits_fcn = 1'h0; // @[top.scala 34:22]
  assign io_imem_req_bits_typ = 3'h7; // @[top.scala 34:22]
  assign assert_out = core__GEN_463;
  assign auto_cover_out = {_GEN_1232,profilePin_615};
  assign core_clock = clock;
  assign core_reset = reset; // @[top.scala 44:28]
  assign core_io_imem_resp_bits_data = io_imem_resp_bits_data; // @[top.scala 34:22]
  assign core_io_dmem_resp_bits_data = memory_io_core_ports_0_resp_bits_data; // @[top.scala 33:22]
  assign memory_clock = clock;
  assign memory_io_core_ports_0_req_bits_addr = core_io_dmem_req_bits_addr; // @[top.scala 33:22]
  assign memory_io_core_ports_0_req_bits_data = core_io_dmem_req_bits_data; // @[top.scala 33:22]
  assign memory_io_core_ports_0_req_bits_fcn = core_io_dmem_req_bits_fcn; // @[top.scala 33:22]
  assign memory_io_core_ports_0_req_bits_typ = core_io_dmem_req_bits_typ; // @[top.scala 33:22]
endmodule
module FrontEnd(
  input         metaReset,
  input         clock,
  input         reset,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_pc,
  input         io_cpu_resp_ready,
  output        io_cpu_resp_valid,
  output [31:0] io_cpu_resp_bits_pc,
  output [31:0] io_cpu_resp_bits_inst,
  output [31:0] io_imem_req_bits_addr,
  input  [31:0] io_imem_resp_bits_data,
  output        _GEN_1_1,
  output        _GEN_10_1,
  output        _GEN_13_1,
  output        _GEN_7_1,
  output        _GEN_9_2,
  output        _GEN_12_3,
  output        _GEN_6_3,
  output        _GEN_5_4,
  output        _GEN_8_3,
  output        _GEN_11_4
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg  if_reg_valid; // @[frontend.scala 87:27]
  wire [31:0] _T_132 = 32'h80000000 - 32'h4; // @[frontend.scala 88:45]
  reg [31:0] if_reg_pc; // @[frontend.scala 88:27]
  reg  exe_reg_valid; // @[frontend.scala 90:27]
  reg [31:0] exe_reg_pc; // @[frontend.scala 91:27]
  reg [31:0] exe_reg_inst; // @[frontend.scala 92:27]
  wire [31:0] if_pc_plus4 = if_reg_pc + 32'h4; // @[frontend.scala 100:33]
  wire [31:0] _GEN_0 = io_cpu_req_valid ? io_cpu_req_bits_pc : if_pc_plus4; // @[frontend.scala 107:7]
  wire  _GEN_3 = io_cpu_resp_ready | if_reg_valid; // @[frontend.scala 118:4]
  wire  _T_144 = ~io_cpu_req_valid; // @[frontend.scala 133:40]
  wire  _T_145 = if_reg_valid & _T_144; // @[frontend.scala 133:37]
  assign io_cpu_resp_valid = exe_reg_valid; // @[frontend.scala 141:26]
  assign io_cpu_resp_bits_pc = exe_reg_pc; // @[frontend.scala 143:26]
  assign io_cpu_resp_bits_inst = exe_reg_inst; // @[frontend.scala 142:26]
  assign io_imem_req_bits_addr = io_cpu_resp_ready ? _GEN_0 : if_reg_pc; // @[frontend.scala 124:26]
  assign _GEN_1_1 = io_cpu_req_valid;
  assign _GEN_10_1 = reset;
  assign _GEN_13_1 = io_cpu_resp_ready;
  assign _GEN_7_1 = io_cpu_resp_ready;
  assign _GEN_9_2 = reset;
  assign _GEN_12_3 = io_cpu_resp_ready;
  assign _GEN_6_3 = io_cpu_resp_ready;
  assign _GEN_5_4 = io_cpu_resp_ready;
  assign _GEN_8_3 = io_cpu_resp_ready;
  assign _GEN_11_4 = reset;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  if_reg_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  if_reg_pc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  exe_reg_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  exe_reg_pc = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  exe_reg_inst = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      if_reg_valid <= 1'h0;
    end else if (reset) begin
      if_reg_valid <= 1'h0;
    end else begin
      if_reg_valid <= _GEN_3;
    end
    if (metaReset) begin
      if_reg_pc <= 32'h0;
    end else if (reset) begin
      if_reg_pc <= _T_132;
    end else if (io_cpu_resp_ready) begin
      if (io_cpu_resp_ready) begin
        if (io_cpu_req_valid) begin
          if_reg_pc <= io_cpu_req_bits_pc;
        end else begin
          if_reg_pc <= if_pc_plus4;
        end
      end
    end
    if (metaReset) begin
      exe_reg_valid <= 1'h0;
    end else if (reset) begin
      exe_reg_valid <= 1'h0;
    end else if (io_cpu_resp_ready) begin
      exe_reg_valid <= _T_145;
    end
    if (metaReset) begin
      exe_reg_pc <= 32'h0;
    end else if (io_cpu_resp_ready) begin
      exe_reg_pc <= if_reg_pc;
    end
    if (metaReset) begin
      exe_reg_inst <= 32'h0;
    end else if (io_cpu_resp_ready) begin
      exe_reg_inst <= io_imem_resp_bits_data;
    end
  end
endmodule
module CtlPath(
  input         metaReset,
  input         clock,
  output        io_imem_req_valid,
  input         io_imem_resp_valid,
  input  [31:0] io_imem_resp_bits_inst,
  input         io_dat_br_eq,
  input         io_dat_br_lt,
  input         io_dat_br_ltu,
  input         io_dat_csr_eret,
  output        io_ctl_exe_kill,
  output [2:0]  io_ctl_pc_sel,
  output        io_ctl_brjmp_sel,
  output [1:0]  io_ctl_op1_sel,
  output [1:0]  io_ctl_op2_sel,
  output [3:0]  io_ctl_alu_fun,
  output [1:0]  io_ctl_wb_sel,
  output        io_ctl_rf_wen,
  output        io_ctl_bypassable,
  output [2:0]  io_ctl_csr_cmd,
  output        io_ctl_dmem_fcn,
  output [2:0]  io_ctl_dmem_typ,
  output        io_ctl_exception,
  output        _GEN_92_0,
  output        _GEN_52_0,
  output        _GEN_305_0,
  output        _GEN_200_0,
  output        _GEN_149_0,
  output        _GEN_25_0,
  output        _GEN_248_0,
  output        _GEN_107_0,
  output        _GEN_134_0,
  output        _GEN_206_0,
  output        _GEN_40_0,
  output        _GEN_233_0,
  output        _GEN_128_0,
  output        _GEN_191_0,
  output        _GEN_227_0,
  output        _GEN_113_0,
  output        _GEN_46_0,
  output        _GEN_299_0,
  output        _GEN_73_0,
  output        _GEN_212_0,
  output        _GEN_31_0,
  output        _GEN_311_0,
  output        _GEN_67_0,
  output        _GEN_320_0,
  output        _GEN_215_0,
  output        _GEN_221_0,
  output        _GEN_101_0,
  output        _GEN_110_0,
  output        _GEN_283_0,
  output        _GEN_314_0,
  output        _GEN_178_0,
  output        _GEN_209_0,
  output        _GEN_28_0,
  output        _GEN_277_0,
  output        _GEN_55_0,
  output        _GEN_194_0,
  output        _GEN_13_0,
  output        _GEN_49_0,
  output        _GEN_116_0,
  output        _GEN_7_0,
  output        _GEN_34_0,
  output        _GEN_122_0,
  output        _GEN_308_0,
  output        _GEN_95_0,
  output        _GEN_230_0,
  output        _GEN_293_0,
  output        _GEN_184_0,
  output        _GEN_1_2,
  output        _GEN_197_0,
  output        _GEN_187_0,
  output        _GEN_104_0,
  output        _GEN_265_0,
  output        _GEN_296_0,
  output        _GEN_160_0,
  output        _GEN_172_0,
  output        _GEN_203_0,
  output        _GEN_271_0,
  output        _GEN_37_0,
  output        _GEN_166_0,
  output        _GEN_280_0,
  output        _GEN_286_0,
  output        _GEN_22_1,
  output        _GEN_302_0,
  output        _GEN_16_2,
  output        _GEN_10_2,
  output        _GEN_259_0,
  output        _GEN_98_0,
  output        _GEN_19_1,
  output        _GEN_148_0,
  output        _GEN_87_0,
  output        _GEN_274_0,
  output        _GEN_232_0,
  output        _GEN_190_0,
  output        _GEN_154_0,
  output        _GEN_289_0,
  output        _GEN_181_0,
  output        _GEN_253_0,
  output        _GEN_72_0,
  output        _GEN_175_0,
  output        _GEN_169_0,
  output        _GEN_4_1,
  output        _GEN_247_0,
  output        _GEN_268_0,
  output        _GEN_214_0,
  output        _GEN_250_0,
  output        _GEN_241_0,
  output        _GEN_142_0,
  output        _GEN_136_0,
  output        _GEN_235_0,
  output        _GEN_262_0,
  output        _GEN_54_0,
  output        _GEN_313_0,
  output        _GEN_69_0,
  output        _GEN_157_0,
  output        _GEN_75_0,
  output        _GEN_90_0,
  output        _GEN_163_0,
  output        _GEN_130_0,
  output        _GEN_229_0,
  output        _GEN_121_0,
  output        _GEN_256_0,
  output        _GEN_81_0,
  output        _GEN_57_0,
  output        _GEN_145_0,
  output        _GEN_223_0,
  output        _GEN_118_0,
  output        _GEN_322_0,
  output        _GEN_244_0,
  output        _GEN_124_0,
  output        _GEN_103_0,
  output        _GEN_238_0,
  output        _GEN_63_0,
  output        _GEN_151_0,
  output        _GEN_202_0,
  output        _GEN_196_0,
  output        _GEN_295_0,
  output        _GEN_301_0,
  output        _GEN_310_0,
  output        _GEN_78_0,
  output        _GEN_84_0,
  output        _GEN_217_0,
  output        _GEN_36_0,
  output        _GEN_42_0,
  output        _GEN_316_0,
  output        _GEN_139_0,
  output        _GEN_18_1,
  output        _GEN_226_0,
  output        _GEN_106_0,
  output        _GEN_51_0,
  output        _GEN_45_0,
  output        _GEN_319_0,
  output        _GEN_39_0,
  output        _GEN_66_0,
  output        _GEN_24_0,
  output        _GEN_112_0,
  output        _GEN_211_0,
  output        _GEN_220_0,
  output        _GEN_133_0,
  output        _GEN_127_0,
  output        _GEN_288_1,
  output        _GEN_91_0,
  output        _GEN_205_0,
  output        _GEN_100_0,
  output        _GEN_304_0,
  output        _GEN_60_0,
  output        _GEN_298_0,
  output        _GEN_189_0,
  output        _GEN_199_0,
  output        _GEN_177_0,
  output        _GEN_12_2,
  output        _GEN_94_0,
  output        _GEN_162_0,
  output        _GEN_193_0,
  output        _GEN_208_0,
  output        _GEN_261_0,
  output        _GEN_115_0,
  output        _GEN_27_0,
  output        _GEN_270_0,
  output        _GEN_183_0,
  output        _GEN_33_0,
  output        _GEN_276_0,
  output        _GEN_282_1,
  output        _GEN_292_0,
  output        _GEN_48_0,
  output        _GEN_6_2,
  output        _GEN_307_0,
  output        _GEN_109_0,
  output        _GEN_21_1,
  output        _GEN_15_3,
  output        _GEN_30_0,
  output        _GEN_83_0,
  output        _GEN_171_0,
  output        _GEN_186_0,
  output        _GEN_144_0,
  output        _GEN_279_1,
  output        _GEN_97_0,
  output        _GEN_264_0,
  output        _GEN_165_0,
  output        _GEN_159_0,
  output        _GEN_258_0,
  output        _GEN_285_1,
  output        _GEN_180_0,
  output        _GEN_9_3,
  output        _GEN_243_0,
  output        _GEN_77_0,
  output        _GEN_174_0,
  output        _GEN_225_0,
  output        _GEN_252_0,
  output        _GEN_132_0,
  output        _GEN_147_1,
  output        _GEN_240_0,
  output        _GEN_65_0,
  output        _GEN_273_0,
  output        _GEN_59_0,
  output        _GEN_231_0,
  output        _GEN_86_0,
  output        _GEN_80_0,
  output        _GEN_3_2,
  output        _GEN_246_0,
  output        _GEN_71_0,
  output        _GEN_153_0,
  output        _GEN_168_0,
  output        _GEN_267_0,
  output        _GEN_126_0,
  output        _GEN_213_0,
  output        _GEN_255_0,
  output        _GEN_156_0,
  output        _GEN_150_0,
  output        _GEN_114_0,
  output        _GEN_228_0,
  output        _GEN_141_0,
  output        _GEN_108_0,
  output        _GEN_249_0,
  output        _GEN_312_1,
  output        _GEN_68_0,
  output        _GEN_74_0,
  output        _GEN_207_0,
  output        _GEN_234_0,
  output        _GEN_306_1,
  output        _GEN_129_0,
  output        _GEN_89_0,
  output        _GEN_47_0,
  output        _GEN_53_0,
  output        _GEN_135_0,
  output        _GEN_222_0,
  output        _GEN_29_0,
  output        _GEN_41_0,
  output        _GEN_56_0,
  output        _GEN_195_0,
  output        _GEN_237_0,
  output        _GEN_102_0,
  output        _GEN_62_0,
  output        _GEN_35_0,
  output        _GEN_123_0,
  output        _GEN_117_0,
  output        _GEN_321_0,
  output        _GEN_216_0,
  output        _GEN_294_1,
  output        _GEN_50_0,
  output        _GEN_138_0,
  output        _GEN_201_0,
  output        _GEN_210_0,
  output        _GEN_96_0,
  output        _GEN_315_0,
  output        _GEN_309_0,
  output        _GEN_17_1,
  output        _GEN_105_0,
  output        _GEN_303_0,
  output        _GEN_204_0,
  output        _GEN_318_1,
  output        _GEN_173_0,
  output        _GEN_198_0,
  output        _GEN_23_1,
  output        _GEN_272_1,
  output        _GEN_120_0,
  output        _GEN_188_0,
  output        _GEN_44_0,
  output        _GEN_287_1,
  output        _GEN_297_0,
  output        _GEN_2_2,
  output        _GEN_99_0,
  output        _GEN_38_0,
  output        _GEN_111_0,
  output        _GEN_219_0,
  output        _GEN_26_0,
  output        _GEN_176_0,
  output        _GEN_182_0,
  output        _GEN_290_1,
  output        _GEN_0_2,
  output        _GEN_32_0,
  output        _GEN_161_0,
  output        _GEN_275_1,
  output        _GEN_170_0,
  output        _GEN_192_0,
  output        _GEN_20_1,
  output        _GEN_269_1,
  output        _GEN_281_1,
  output        _GEN_291_1,
  output        _GEN_155_0,
  output        _GEN_88_0,
  output        _GEN_300_1,
  output        _GEN_11_3,
  output        _GEN_5_3,
  output        _GEN_254_1,
  output        _GEN_93_0,
  output        _GEN_14_2,
  output        _GEN_257_1,
  output        _GEN_82_0,
  output        _GEN_8_2,
  output        _GEN_278_1,
  output        _GEN_70_0,
  output        _GEN_158_0,
  output        _GEN_236_1,
  output        _GEN_185_0,
  output        _GEN_61_0,
  output        _GEN_143_0,
  output        _GEN_284_1,
  output        _GEN_179_0,
  output        _GEN_242_1,
  output        _GEN_137_0,
  output        _GEN_76_0,
  output        _GEN_164_0,
  output        _GEN_263_1,
  output        _GEN_167_0,
  output        _GEN_43_0,
  output        _GEN_266_1,
  output        _GEN_131_0,
  output        _GEN_125_0,
  output        _GEN_317_1,
  output        _GEN_224_0,
  output        _GEN_119_0,
  output        _GEN_239_1,
  output        _GEN_152_1,
  output        _GEN_146_1,
  output        _GEN_245_1,
  output        _GEN_323_1,
  output        _GEN_79_0,
  output        _GEN_218_0,
  output        _GEN_64_0,
  output        _GEN_58_0,
  output        _GEN_251_1,
  output        _GEN_260_1,
  output        _GEN_140_0,
  output        _GEN_85_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] _T_88 = io_imem_resp_bits_inst & 32'h707f; // @[Lookup.scala 9:38]
  wire  _T_89 = 32'h2003 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_93 = 32'h3 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_97 = 32'h4003 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_101 = 32'h1003 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_105 = 32'h5003 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_109 = 32'h2023 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_113 = 32'h23 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_117 = 32'h1023 == _T_88; // @[Lookup.scala 9:38]
  wire [31:0] _T_120 = io_imem_resp_bits_inst & 32'h7f; // @[Lookup.scala 9:38]
  wire  _T_121 = 32'h17 == _T_120; // @[Lookup.scala 9:38]
  wire  _T_125 = 32'h37 == _T_120; // @[Lookup.scala 9:38]
  wire  _T_129 = 32'h13 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_133 = 32'h7013 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_137 = 32'h6013 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_141 = 32'h4013 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_145 = 32'h2013 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_149 = 32'h3013 == _T_88; // @[Lookup.scala 9:38]
  wire [31:0] _T_152 = io_imem_resp_bits_inst & 32'hfc00707f; // @[Lookup.scala 9:38]
  wire  _T_153 = 32'h1013 == _T_152; // @[Lookup.scala 9:38]
  wire  _T_157 = 32'h40005013 == _T_152; // @[Lookup.scala 9:38]
  wire  _T_161 = 32'h5013 == _T_152; // @[Lookup.scala 9:38]
  wire [31:0] _T_164 = io_imem_resp_bits_inst & 32'hfe00707f; // @[Lookup.scala 9:38]
  wire  _T_165 = 32'h1033 == _T_164; // @[Lookup.scala 9:38]
  wire  _T_169 = 32'h33 == _T_164; // @[Lookup.scala 9:38]
  wire  _T_173 = 32'h40000033 == _T_164; // @[Lookup.scala 9:38]
  wire  _T_177 = 32'h2033 == _T_164; // @[Lookup.scala 9:38]
  wire  _T_181 = 32'h3033 == _T_164; // @[Lookup.scala 9:38]
  wire  _T_185 = 32'h7033 == _T_164; // @[Lookup.scala 9:38]
  wire  _T_189 = 32'h6033 == _T_164; // @[Lookup.scala 9:38]
  wire  _T_193 = 32'h4033 == _T_164; // @[Lookup.scala 9:38]
  wire  _T_197 = 32'h40005033 == _T_164; // @[Lookup.scala 9:38]
  wire  _T_201 = 32'h5033 == _T_164; // @[Lookup.scala 9:38]
  wire  _T_205 = 32'h6f == _T_120; // @[Lookup.scala 9:38]
  wire  _T_209 = 32'h67 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_213 = 32'h63 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_217 = 32'h1063 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_221 = 32'h5063 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_225 = 32'h7063 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_229 = 32'h4063 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_233 = 32'h6063 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_237 = 32'h5073 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_241 = 32'h6073 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_245 = 32'h1073 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_249 = 32'h2073 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_253 = 32'h3073 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_257 = 32'h7073 == _T_88; // @[Lookup.scala 9:38]
  wire  _T_261 = 32'h73 == io_imem_resp_bits_inst; // @[Lookup.scala 9:38]
  wire  _T_265 = 32'h30200073 == io_imem_resp_bits_inst; // @[Lookup.scala 9:38]
  wire  _T_269 = 32'h7b200073 == io_imem_resp_bits_inst; // @[Lookup.scala 9:38]
  wire  _T_273 = 32'h100073 == io_imem_resp_bits_inst; // @[Lookup.scala 9:38]
  wire  _T_277 = 32'h10500073 == io_imem_resp_bits_inst; // @[Lookup.scala 9:38]
  wire  _T_281 = 32'h100f == _T_88; // @[Lookup.scala 9:38]
  wire  _T_285 = 32'hf == _T_88; // @[Lookup.scala 9:38]
  wire  _T_287 = _T_281 | _T_285; // @[Lookup.scala 11:37]
  wire  _T_288 = _T_277 | _T_287; // @[Lookup.scala 11:37]
  wire  _T_289 = _T_273 | _T_288; // @[Lookup.scala 11:37]
  wire  _T_290 = _T_269 | _T_289; // @[Lookup.scala 11:37]
  wire  _T_291 = _T_265 | _T_290; // @[Lookup.scala 11:37]
  wire  _T_292 = _T_261 | _T_291; // @[Lookup.scala 11:37]
  wire  _T_293 = _T_257 | _T_292; // @[Lookup.scala 11:37]
  wire  _T_294 = _T_253 | _T_293; // @[Lookup.scala 11:37]
  wire  _T_295 = _T_249 | _T_294; // @[Lookup.scala 11:37]
  wire  _T_296 = _T_245 | _T_295; // @[Lookup.scala 11:37]
  wire  _T_297 = _T_241 | _T_296; // @[Lookup.scala 11:37]
  wire  _T_298 = _T_237 | _T_297; // @[Lookup.scala 11:37]
  wire  _T_299 = _T_233 | _T_298; // @[Lookup.scala 11:37]
  wire  _T_300 = _T_229 | _T_299; // @[Lookup.scala 11:37]
  wire  _T_301 = _T_225 | _T_300; // @[Lookup.scala 11:37]
  wire  _T_302 = _T_221 | _T_301; // @[Lookup.scala 11:37]
  wire  _T_303 = _T_217 | _T_302; // @[Lookup.scala 11:37]
  wire  _T_304 = _T_213 | _T_303; // @[Lookup.scala 11:37]
  wire  _T_305 = _T_209 | _T_304; // @[Lookup.scala 11:37]
  wire  _T_306 = _T_205 | _T_305; // @[Lookup.scala 11:37]
  wire  _T_307 = _T_201 | _T_306; // @[Lookup.scala 11:37]
  wire  _T_308 = _T_197 | _T_307; // @[Lookup.scala 11:37]
  wire  _T_309 = _T_193 | _T_308; // @[Lookup.scala 11:37]
  wire  _T_310 = _T_189 | _T_309; // @[Lookup.scala 11:37]
  wire  _T_311 = _T_185 | _T_310; // @[Lookup.scala 11:37]
  wire  _T_312 = _T_181 | _T_311; // @[Lookup.scala 11:37]
  wire  _T_313 = _T_177 | _T_312; // @[Lookup.scala 11:37]
  wire  _T_314 = _T_173 | _T_313; // @[Lookup.scala 11:37]
  wire  _T_315 = _T_169 | _T_314; // @[Lookup.scala 11:37]
  wire  _T_316 = _T_165 | _T_315; // @[Lookup.scala 11:37]
  wire  _T_317 = _T_161 | _T_316; // @[Lookup.scala 11:37]
  wire  _T_318 = _T_157 | _T_317; // @[Lookup.scala 11:37]
  wire  _T_319 = _T_153 | _T_318; // @[Lookup.scala 11:37]
  wire  _T_320 = _T_149 | _T_319; // @[Lookup.scala 11:37]
  wire  _T_321 = _T_145 | _T_320; // @[Lookup.scala 11:37]
  wire  _T_322 = _T_141 | _T_321; // @[Lookup.scala 11:37]
  wire  _T_323 = _T_137 | _T_322; // @[Lookup.scala 11:37]
  wire  _T_324 = _T_133 | _T_323; // @[Lookup.scala 11:37]
  wire  _T_325 = _T_129 | _T_324; // @[Lookup.scala 11:37]
  wire  _T_326 = _T_125 | _T_325; // @[Lookup.scala 11:37]
  wire  _T_327 = _T_121 | _T_326; // @[Lookup.scala 11:37]
  wire  _T_328 = _T_117 | _T_327; // @[Lookup.scala 11:37]
  wire  _T_329 = _T_113 | _T_328; // @[Lookup.scala 11:37]
  wire  _T_330 = _T_109 | _T_329; // @[Lookup.scala 11:37]
  wire  _T_331 = _T_105 | _T_330; // @[Lookup.scala 11:37]
  wire  _T_332 = _T_101 | _T_331; // @[Lookup.scala 11:37]
  wire  _T_333 = _T_97 | _T_332; // @[Lookup.scala 11:37]
  wire  _T_334 = _T_93 | _T_333; // @[Lookup.scala 11:37]
  wire  cs_inst_val = _T_89 | _T_334; // @[Lookup.scala 11:37]
  wire [3:0] _T_348 = _T_233 ? 4'h6 : 4'h0; // @[Lookup.scala 11:37]
  wire [3:0] _T_349 = _T_229 ? 4'h5 : _T_348; // @[Lookup.scala 11:37]
  wire [3:0] _T_350 = _T_225 ? 4'h4 : _T_349; // @[Lookup.scala 11:37]
  wire [3:0] _T_351 = _T_221 ? 4'h3 : _T_350; // @[Lookup.scala 11:37]
  wire [3:0] _T_352 = _T_217 ? 4'h1 : _T_351; // @[Lookup.scala 11:37]
  wire [3:0] _T_353 = _T_213 ? 4'h2 : _T_352; // @[Lookup.scala 11:37]
  wire [3:0] _T_354 = _T_209 ? 4'h8 : _T_353; // @[Lookup.scala 11:37]
  wire [3:0] _T_355 = _T_205 ? 4'h7 : _T_354; // @[Lookup.scala 11:37]
  wire [3:0] _T_356 = _T_201 ? 4'h0 : _T_355; // @[Lookup.scala 11:37]
  wire [3:0] _T_357 = _T_197 ? 4'h0 : _T_356; // @[Lookup.scala 11:37]
  wire [3:0] _T_358 = _T_193 ? 4'h0 : _T_357; // @[Lookup.scala 11:37]
  wire [3:0] _T_359 = _T_189 ? 4'h0 : _T_358; // @[Lookup.scala 11:37]
  wire [3:0] _T_360 = _T_185 ? 4'h0 : _T_359; // @[Lookup.scala 11:37]
  wire [3:0] _T_361 = _T_181 ? 4'h0 : _T_360; // @[Lookup.scala 11:37]
  wire [3:0] _T_362 = _T_177 ? 4'h0 : _T_361; // @[Lookup.scala 11:37]
  wire [3:0] _T_363 = _T_173 ? 4'h0 : _T_362; // @[Lookup.scala 11:37]
  wire [3:0] _T_364 = _T_169 ? 4'h0 : _T_363; // @[Lookup.scala 11:37]
  wire [3:0] _T_365 = _T_165 ? 4'h0 : _T_364; // @[Lookup.scala 11:37]
  wire [3:0] _T_366 = _T_161 ? 4'h0 : _T_365; // @[Lookup.scala 11:37]
  wire [3:0] _T_367 = _T_157 ? 4'h0 : _T_366; // @[Lookup.scala 11:37]
  wire [3:0] _T_368 = _T_153 ? 4'h0 : _T_367; // @[Lookup.scala 11:37]
  wire [3:0] _T_369 = _T_149 ? 4'h0 : _T_368; // @[Lookup.scala 11:37]
  wire [3:0] _T_370 = _T_145 ? 4'h0 : _T_369; // @[Lookup.scala 11:37]
  wire [3:0] _T_371 = _T_141 ? 4'h0 : _T_370; // @[Lookup.scala 11:37]
  wire [3:0] _T_372 = _T_137 ? 4'h0 : _T_371; // @[Lookup.scala 11:37]
  wire [3:0] _T_373 = _T_133 ? 4'h0 : _T_372; // @[Lookup.scala 11:37]
  wire [3:0] _T_374 = _T_129 ? 4'h0 : _T_373; // @[Lookup.scala 11:37]
  wire [3:0] _T_375 = _T_125 ? 4'h0 : _T_374; // @[Lookup.scala 11:37]
  wire [3:0] _T_376 = _T_121 ? 4'h0 : _T_375; // @[Lookup.scala 11:37]
  wire [3:0] _T_377 = _T_117 ? 4'h0 : _T_376; // @[Lookup.scala 11:37]
  wire [3:0] _T_378 = _T_113 ? 4'h0 : _T_377; // @[Lookup.scala 11:37]
  wire [3:0] _T_379 = _T_109 ? 4'h0 : _T_378; // @[Lookup.scala 11:37]
  wire [3:0] _T_380 = _T_105 ? 4'h0 : _T_379; // @[Lookup.scala 11:37]
  wire [3:0] _T_381 = _T_101 ? 4'h0 : _T_380; // @[Lookup.scala 11:37]
  wire [3:0] _T_382 = _T_97 ? 4'h0 : _T_381; // @[Lookup.scala 11:37]
  wire [3:0] _T_383 = _T_93 ? 4'h0 : _T_382; // @[Lookup.scala 11:37]
  wire [3:0] cs_br_type = _T_89 ? 4'h0 : _T_383; // @[Lookup.scala 11:37]
  wire  _T_404 = _T_205 | _T_209; // @[Lookup.scala 11:37]
  wire  _T_405 = _T_201 ? 1'h0 : _T_404; // @[Lookup.scala 11:37]
  wire  _T_406 = _T_197 ? 1'h0 : _T_405; // @[Lookup.scala 11:37]
  wire  _T_407 = _T_193 ? 1'h0 : _T_406; // @[Lookup.scala 11:37]
  wire  _T_408 = _T_189 ? 1'h0 : _T_407; // @[Lookup.scala 11:37]
  wire  _T_409 = _T_185 ? 1'h0 : _T_408; // @[Lookup.scala 11:37]
  wire  _T_410 = _T_181 ? 1'h0 : _T_409; // @[Lookup.scala 11:37]
  wire  _T_411 = _T_177 ? 1'h0 : _T_410; // @[Lookup.scala 11:37]
  wire  _T_412 = _T_173 ? 1'h0 : _T_411; // @[Lookup.scala 11:37]
  wire  _T_413 = _T_169 ? 1'h0 : _T_412; // @[Lookup.scala 11:37]
  wire  _T_414 = _T_165 ? 1'h0 : _T_413; // @[Lookup.scala 11:37]
  wire  _T_415 = _T_161 ? 1'h0 : _T_414; // @[Lookup.scala 11:37]
  wire  _T_416 = _T_157 ? 1'h0 : _T_415; // @[Lookup.scala 11:37]
  wire  _T_417 = _T_153 ? 1'h0 : _T_416; // @[Lookup.scala 11:37]
  wire  _T_418 = _T_149 ? 1'h0 : _T_417; // @[Lookup.scala 11:37]
  wire  _T_419 = _T_145 ? 1'h0 : _T_418; // @[Lookup.scala 11:37]
  wire  _T_420 = _T_141 ? 1'h0 : _T_419; // @[Lookup.scala 11:37]
  wire  _T_421 = _T_137 ? 1'h0 : _T_420; // @[Lookup.scala 11:37]
  wire  _T_422 = _T_133 ? 1'h0 : _T_421; // @[Lookup.scala 11:37]
  wire  _T_423 = _T_129 ? 1'h0 : _T_422; // @[Lookup.scala 11:37]
  wire  _T_424 = _T_125 ? 1'h0 : _T_423; // @[Lookup.scala 11:37]
  wire  _T_425 = _T_121 ? 1'h0 : _T_424; // @[Lookup.scala 11:37]
  wire  _T_426 = _T_117 ? 1'h0 : _T_425; // @[Lookup.scala 11:37]
  wire  _T_427 = _T_113 ? 1'h0 : _T_426; // @[Lookup.scala 11:37]
  wire  _T_428 = _T_109 ? 1'h0 : _T_427; // @[Lookup.scala 11:37]
  wire  _T_429 = _T_105 ? 1'h0 : _T_428; // @[Lookup.scala 11:37]
  wire  _T_430 = _T_101 ? 1'h0 : _T_429; // @[Lookup.scala 11:37]
  wire  _T_431 = _T_97 ? 1'h0 : _T_430; // @[Lookup.scala 11:37]
  wire  _T_432 = _T_93 ? 1'h0 : _T_431; // @[Lookup.scala 11:37]
  wire [1:0] _T_440 = _T_257 ? 2'h2 : 2'h0; // @[Lookup.scala 11:37]
  wire [1:0] _T_441 = _T_253 ? 2'h0 : _T_440; // @[Lookup.scala 11:37]
  wire [1:0] _T_442 = _T_249 ? 2'h0 : _T_441; // @[Lookup.scala 11:37]
  wire [1:0] _T_443 = _T_245 ? 2'h0 : _T_442; // @[Lookup.scala 11:37]
  wire [1:0] _T_444 = _T_241 ? 2'h2 : _T_443; // @[Lookup.scala 11:37]
  wire [1:0] _T_445 = _T_237 ? 2'h2 : _T_444; // @[Lookup.scala 11:37]
  wire [1:0] _T_446 = _T_233 ? 2'h0 : _T_445; // @[Lookup.scala 11:37]
  wire [1:0] _T_447 = _T_229 ? 2'h0 : _T_446; // @[Lookup.scala 11:37]
  wire [1:0] _T_448 = _T_225 ? 2'h0 : _T_447; // @[Lookup.scala 11:37]
  wire [1:0] _T_449 = _T_221 ? 2'h0 : _T_448; // @[Lookup.scala 11:37]
  wire [1:0] _T_450 = _T_217 ? 2'h0 : _T_449; // @[Lookup.scala 11:37]
  wire [1:0] _T_451 = _T_213 ? 2'h0 : _T_450; // @[Lookup.scala 11:37]
  wire [1:0] _T_452 = _T_209 ? 2'h0 : _T_451; // @[Lookup.scala 11:37]
  wire [1:0] _T_453 = _T_205 ? 2'h0 : _T_452; // @[Lookup.scala 11:37]
  wire [1:0] _T_454 = _T_201 ? 2'h0 : _T_453; // @[Lookup.scala 11:37]
  wire [1:0] _T_455 = _T_197 ? 2'h0 : _T_454; // @[Lookup.scala 11:37]
  wire [1:0] _T_456 = _T_193 ? 2'h0 : _T_455; // @[Lookup.scala 11:37]
  wire [1:0] _T_457 = _T_189 ? 2'h0 : _T_456; // @[Lookup.scala 11:37]
  wire [1:0] _T_458 = _T_185 ? 2'h0 : _T_457; // @[Lookup.scala 11:37]
  wire [1:0] _T_459 = _T_181 ? 2'h0 : _T_458; // @[Lookup.scala 11:37]
  wire [1:0] _T_460 = _T_177 ? 2'h0 : _T_459; // @[Lookup.scala 11:37]
  wire [1:0] _T_461 = _T_173 ? 2'h0 : _T_460; // @[Lookup.scala 11:37]
  wire [1:0] _T_462 = _T_169 ? 2'h0 : _T_461; // @[Lookup.scala 11:37]
  wire [1:0] _T_463 = _T_165 ? 2'h0 : _T_462; // @[Lookup.scala 11:37]
  wire [1:0] _T_464 = _T_161 ? 2'h0 : _T_463; // @[Lookup.scala 11:37]
  wire [1:0] _T_465 = _T_157 ? 2'h0 : _T_464; // @[Lookup.scala 11:37]
  wire [1:0] _T_466 = _T_153 ? 2'h0 : _T_465; // @[Lookup.scala 11:37]
  wire [1:0] _T_467 = _T_149 ? 2'h0 : _T_466; // @[Lookup.scala 11:37]
  wire [1:0] _T_468 = _T_145 ? 2'h0 : _T_467; // @[Lookup.scala 11:37]
  wire [1:0] _T_469 = _T_141 ? 2'h0 : _T_468; // @[Lookup.scala 11:37]
  wire [1:0] _T_470 = _T_137 ? 2'h0 : _T_469; // @[Lookup.scala 11:37]
  wire [1:0] _T_471 = _T_133 ? 2'h0 : _T_470; // @[Lookup.scala 11:37]
  wire [1:0] _T_472 = _T_129 ? 2'h0 : _T_471; // @[Lookup.scala 11:37]
  wire [1:0] _T_473 = _T_125 ? 2'h1 : _T_472; // @[Lookup.scala 11:37]
  wire [1:0] _T_474 = _T_121 ? 2'h1 : _T_473; // @[Lookup.scala 11:37]
  wire [1:0] _T_475 = _T_117 ? 2'h0 : _T_474; // @[Lookup.scala 11:37]
  wire [1:0] _T_476 = _T_113 ? 2'h0 : _T_475; // @[Lookup.scala 11:37]
  wire [1:0] _T_477 = _T_109 ? 2'h0 : _T_476; // @[Lookup.scala 11:37]
  wire [1:0] _T_478 = _T_105 ? 2'h0 : _T_477; // @[Lookup.scala 11:37]
  wire [1:0] _T_479 = _T_101 ? 2'h0 : _T_478; // @[Lookup.scala 11:37]
  wire [1:0] _T_480 = _T_97 ? 2'h0 : _T_479; // @[Lookup.scala 11:37]
  wire [1:0] _T_481 = _T_93 ? 2'h0 : _T_480; // @[Lookup.scala 11:37]
  wire [1:0] _T_501 = _T_209 ? 2'h1 : 2'h0; // @[Lookup.scala 11:37]
  wire [1:0] _T_502 = _T_205 ? 2'h0 : _T_501; // @[Lookup.scala 11:37]
  wire [1:0] _T_503 = _T_201 ? 2'h0 : _T_502; // @[Lookup.scala 11:37]
  wire [1:0] _T_504 = _T_197 ? 2'h0 : _T_503; // @[Lookup.scala 11:37]
  wire [1:0] _T_505 = _T_193 ? 2'h0 : _T_504; // @[Lookup.scala 11:37]
  wire [1:0] _T_506 = _T_189 ? 2'h0 : _T_505; // @[Lookup.scala 11:37]
  wire [1:0] _T_507 = _T_185 ? 2'h0 : _T_506; // @[Lookup.scala 11:37]
  wire [1:0] _T_508 = _T_181 ? 2'h0 : _T_507; // @[Lookup.scala 11:37]
  wire [1:0] _T_509 = _T_177 ? 2'h0 : _T_508; // @[Lookup.scala 11:37]
  wire [1:0] _T_510 = _T_173 ? 2'h0 : _T_509; // @[Lookup.scala 11:37]
  wire [1:0] _T_511 = _T_169 ? 2'h0 : _T_510; // @[Lookup.scala 11:37]
  wire [1:0] _T_512 = _T_165 ? 2'h0 : _T_511; // @[Lookup.scala 11:37]
  wire [1:0] _T_513 = _T_161 ? 2'h1 : _T_512; // @[Lookup.scala 11:37]
  wire [1:0] _T_514 = _T_157 ? 2'h1 : _T_513; // @[Lookup.scala 11:37]
  wire [1:0] _T_515 = _T_153 ? 2'h1 : _T_514; // @[Lookup.scala 11:37]
  wire [1:0] _T_516 = _T_149 ? 2'h1 : _T_515; // @[Lookup.scala 11:37]
  wire [1:0] _T_517 = _T_145 ? 2'h1 : _T_516; // @[Lookup.scala 11:37]
  wire [1:0] _T_518 = _T_141 ? 2'h1 : _T_517; // @[Lookup.scala 11:37]
  wire [1:0] _T_519 = _T_137 ? 2'h1 : _T_518; // @[Lookup.scala 11:37]
  wire [1:0] _T_520 = _T_133 ? 2'h1 : _T_519; // @[Lookup.scala 11:37]
  wire [1:0] _T_521 = _T_129 ? 2'h1 : _T_520; // @[Lookup.scala 11:37]
  wire [1:0] _T_522 = _T_125 ? 2'h0 : _T_521; // @[Lookup.scala 11:37]
  wire [1:0] _T_523 = _T_121 ? 2'h3 : _T_522; // @[Lookup.scala 11:37]
  wire [1:0] _T_524 = _T_117 ? 2'h2 : _T_523; // @[Lookup.scala 11:37]
  wire [1:0] _T_525 = _T_113 ? 2'h2 : _T_524; // @[Lookup.scala 11:37]
  wire [1:0] _T_526 = _T_109 ? 2'h2 : _T_525; // @[Lookup.scala 11:37]
  wire [1:0] _T_527 = _T_105 ? 2'h1 : _T_526; // @[Lookup.scala 11:37]
  wire [1:0] _T_528 = _T_101 ? 2'h1 : _T_527; // @[Lookup.scala 11:37]
  wire [1:0] _T_529 = _T_97 ? 2'h1 : _T_528; // @[Lookup.scala 11:37]
  wire [1:0] _T_530 = _T_93 ? 2'h1 : _T_529; // @[Lookup.scala 11:37]
  wire [3:0] _T_538 = _T_257 ? 4'h8 : 4'h0; // @[Lookup.scala 11:37]
  wire [3:0] _T_539 = _T_253 ? 4'h8 : _T_538; // @[Lookup.scala 11:37]
  wire [3:0] _T_540 = _T_249 ? 4'h8 : _T_539; // @[Lookup.scala 11:37]
  wire [3:0] _T_541 = _T_245 ? 4'h8 : _T_540; // @[Lookup.scala 11:37]
  wire [3:0] _T_542 = _T_241 ? 4'h8 : _T_541; // @[Lookup.scala 11:37]
  wire [3:0] _T_543 = _T_237 ? 4'h8 : _T_542; // @[Lookup.scala 11:37]
  wire [3:0] _T_544 = _T_233 ? 4'h0 : _T_543; // @[Lookup.scala 11:37]
  wire [3:0] _T_545 = _T_229 ? 4'h0 : _T_544; // @[Lookup.scala 11:37]
  wire [3:0] _T_546 = _T_225 ? 4'h0 : _T_545; // @[Lookup.scala 11:37]
  wire [3:0] _T_547 = _T_221 ? 4'h0 : _T_546; // @[Lookup.scala 11:37]
  wire [3:0] _T_548 = _T_217 ? 4'h0 : _T_547; // @[Lookup.scala 11:37]
  wire [3:0] _T_549 = _T_213 ? 4'h0 : _T_548; // @[Lookup.scala 11:37]
  wire [3:0] _T_550 = _T_209 ? 4'h0 : _T_549; // @[Lookup.scala 11:37]
  wire [3:0] _T_551 = _T_205 ? 4'h0 : _T_550; // @[Lookup.scala 11:37]
  wire [3:0] _T_552 = _T_201 ? 4'h5 : _T_551; // @[Lookup.scala 11:37]
  wire [3:0] _T_553 = _T_197 ? 4'hb : _T_552; // @[Lookup.scala 11:37]
  wire [3:0] _T_554 = _T_193 ? 4'h4 : _T_553; // @[Lookup.scala 11:37]
  wire [3:0] _T_555 = _T_189 ? 4'h6 : _T_554; // @[Lookup.scala 11:37]
  wire [3:0] _T_556 = _T_185 ? 4'h7 : _T_555; // @[Lookup.scala 11:37]
  wire [3:0] _T_557 = _T_181 ? 4'he : _T_556; // @[Lookup.scala 11:37]
  wire [3:0] _T_558 = _T_177 ? 4'hc : _T_557; // @[Lookup.scala 11:37]
  wire [3:0] _T_559 = _T_173 ? 4'ha : _T_558; // @[Lookup.scala 11:37]
  wire [3:0] _T_560 = _T_169 ? 4'h0 : _T_559; // @[Lookup.scala 11:37]
  wire [3:0] _T_561 = _T_165 ? 4'h1 : _T_560; // @[Lookup.scala 11:37]
  wire [3:0] _T_562 = _T_161 ? 4'h5 : _T_561; // @[Lookup.scala 11:37]
  wire [3:0] _T_563 = _T_157 ? 4'hb : _T_562; // @[Lookup.scala 11:37]
  wire [3:0] _T_564 = _T_153 ? 4'h1 : _T_563; // @[Lookup.scala 11:37]
  wire [3:0] _T_565 = _T_149 ? 4'he : _T_564; // @[Lookup.scala 11:37]
  wire [3:0] _T_566 = _T_145 ? 4'hc : _T_565; // @[Lookup.scala 11:37]
  wire [3:0] _T_567 = _T_141 ? 4'h4 : _T_566; // @[Lookup.scala 11:37]
  wire [3:0] _T_568 = _T_137 ? 4'h6 : _T_567; // @[Lookup.scala 11:37]
  wire [3:0] _T_569 = _T_133 ? 4'h7 : _T_568; // @[Lookup.scala 11:37]
  wire [3:0] _T_570 = _T_129 ? 4'h0 : _T_569; // @[Lookup.scala 11:37]
  wire [3:0] _T_571 = _T_125 ? 4'h8 : _T_570; // @[Lookup.scala 11:37]
  wire [3:0] _T_572 = _T_121 ? 4'h0 : _T_571; // @[Lookup.scala 11:37]
  wire [3:0] _T_573 = _T_117 ? 4'h0 : _T_572; // @[Lookup.scala 11:37]
  wire [3:0] _T_574 = _T_113 ? 4'h0 : _T_573; // @[Lookup.scala 11:37]
  wire [3:0] _T_575 = _T_109 ? 4'h0 : _T_574; // @[Lookup.scala 11:37]
  wire [3:0] _T_576 = _T_105 ? 4'h0 : _T_575; // @[Lookup.scala 11:37]
  wire [3:0] _T_577 = _T_101 ? 4'h0 : _T_576; // @[Lookup.scala 11:37]
  wire [3:0] _T_578 = _T_97 ? 4'h0 : _T_577; // @[Lookup.scala 11:37]
  wire [3:0] _T_579 = _T_93 ? 4'h0 : _T_578; // @[Lookup.scala 11:37]
  wire [1:0] _T_587 = _T_257 ? 2'h3 : 2'h0; // @[Lookup.scala 11:37]
  wire [1:0] _T_588 = _T_253 ? 2'h3 : _T_587; // @[Lookup.scala 11:37]
  wire [1:0] _T_589 = _T_249 ? 2'h3 : _T_588; // @[Lookup.scala 11:37]
  wire [1:0] _T_590 = _T_245 ? 2'h3 : _T_589; // @[Lookup.scala 11:37]
  wire [1:0] _T_591 = _T_241 ? 2'h3 : _T_590; // @[Lookup.scala 11:37]
  wire [1:0] _T_592 = _T_237 ? 2'h3 : _T_591; // @[Lookup.scala 11:37]
  wire [1:0] _T_593 = _T_233 ? 2'h0 : _T_592; // @[Lookup.scala 11:37]
  wire [1:0] _T_594 = _T_229 ? 2'h0 : _T_593; // @[Lookup.scala 11:37]
  wire [1:0] _T_595 = _T_225 ? 2'h0 : _T_594; // @[Lookup.scala 11:37]
  wire [1:0] _T_596 = _T_221 ? 2'h0 : _T_595; // @[Lookup.scala 11:37]
  wire [1:0] _T_597 = _T_217 ? 2'h0 : _T_596; // @[Lookup.scala 11:37]
  wire [1:0] _T_598 = _T_213 ? 2'h0 : _T_597; // @[Lookup.scala 11:37]
  wire [1:0] _T_599 = _T_209 ? 2'h2 : _T_598; // @[Lookup.scala 11:37]
  wire [1:0] _T_600 = _T_205 ? 2'h2 : _T_599; // @[Lookup.scala 11:37]
  wire [1:0] _T_601 = _T_201 ? 2'h0 : _T_600; // @[Lookup.scala 11:37]
  wire [1:0] _T_602 = _T_197 ? 2'h0 : _T_601; // @[Lookup.scala 11:37]
  wire [1:0] _T_603 = _T_193 ? 2'h0 : _T_602; // @[Lookup.scala 11:37]
  wire [1:0] _T_604 = _T_189 ? 2'h0 : _T_603; // @[Lookup.scala 11:37]
  wire [1:0] _T_605 = _T_185 ? 2'h0 : _T_604; // @[Lookup.scala 11:37]
  wire [1:0] _T_606 = _T_181 ? 2'h0 : _T_605; // @[Lookup.scala 11:37]
  wire [1:0] _T_607 = _T_177 ? 2'h0 : _T_606; // @[Lookup.scala 11:37]
  wire [1:0] _T_608 = _T_173 ? 2'h0 : _T_607; // @[Lookup.scala 11:37]
  wire [1:0] _T_609 = _T_169 ? 2'h0 : _T_608; // @[Lookup.scala 11:37]
  wire [1:0] _T_610 = _T_165 ? 2'h0 : _T_609; // @[Lookup.scala 11:37]
  wire [1:0] _T_611 = _T_161 ? 2'h0 : _T_610; // @[Lookup.scala 11:37]
  wire [1:0] _T_612 = _T_157 ? 2'h0 : _T_611; // @[Lookup.scala 11:37]
  wire [1:0] _T_613 = _T_153 ? 2'h0 : _T_612; // @[Lookup.scala 11:37]
  wire [1:0] _T_614 = _T_149 ? 2'h0 : _T_613; // @[Lookup.scala 11:37]
  wire [1:0] _T_615 = _T_145 ? 2'h0 : _T_614; // @[Lookup.scala 11:37]
  wire [1:0] _T_616 = _T_141 ? 2'h0 : _T_615; // @[Lookup.scala 11:37]
  wire [1:0] _T_617 = _T_137 ? 2'h0 : _T_616; // @[Lookup.scala 11:37]
  wire [1:0] _T_618 = _T_133 ? 2'h0 : _T_617; // @[Lookup.scala 11:37]
  wire [1:0] _T_619 = _T_129 ? 2'h0 : _T_618; // @[Lookup.scala 11:37]
  wire [1:0] _T_620 = _T_125 ? 2'h0 : _T_619; // @[Lookup.scala 11:37]
  wire [1:0] _T_621 = _T_121 ? 2'h0 : _T_620; // @[Lookup.scala 11:37]
  wire [1:0] _T_622 = _T_117 ? 2'h0 : _T_621; // @[Lookup.scala 11:37]
  wire [1:0] _T_623 = _T_113 ? 2'h0 : _T_622; // @[Lookup.scala 11:37]
  wire [1:0] _T_624 = _T_109 ? 2'h0 : _T_623; // @[Lookup.scala 11:37]
  wire [1:0] _T_625 = _T_105 ? 2'h1 : _T_624; // @[Lookup.scala 11:37]
  wire [1:0] _T_626 = _T_101 ? 2'h1 : _T_625; // @[Lookup.scala 11:37]
  wire [1:0] _T_627 = _T_97 ? 2'h1 : _T_626; // @[Lookup.scala 11:37]
  wire [1:0] _T_628 = _T_93 ? 2'h1 : _T_627; // @[Lookup.scala 11:37]
  wire  _T_637 = _T_253 | _T_257; // @[Lookup.scala 11:37]
  wire  _T_638 = _T_249 | _T_637; // @[Lookup.scala 11:37]
  wire  _T_639 = _T_245 | _T_638; // @[Lookup.scala 11:37]
  wire  _T_640 = _T_241 | _T_639; // @[Lookup.scala 11:37]
  wire  _T_641 = _T_237 | _T_640; // @[Lookup.scala 11:37]
  wire  _T_642 = _T_233 ? 1'h0 : _T_641; // @[Lookup.scala 11:37]
  wire  _T_643 = _T_229 ? 1'h0 : _T_642; // @[Lookup.scala 11:37]
  wire  _T_644 = _T_225 ? 1'h0 : _T_643; // @[Lookup.scala 11:37]
  wire  _T_645 = _T_221 ? 1'h0 : _T_644; // @[Lookup.scala 11:37]
  wire  _T_646 = _T_217 ? 1'h0 : _T_645; // @[Lookup.scala 11:37]
  wire  _T_647 = _T_213 ? 1'h0 : _T_646; // @[Lookup.scala 11:37]
  wire  _T_648 = _T_209 | _T_647; // @[Lookup.scala 11:37]
  wire  _T_649 = _T_205 | _T_648; // @[Lookup.scala 11:37]
  wire  _T_650 = _T_201 | _T_649; // @[Lookup.scala 11:37]
  wire  _T_651 = _T_197 | _T_650; // @[Lookup.scala 11:37]
  wire  _T_652 = _T_193 | _T_651; // @[Lookup.scala 11:37]
  wire  _T_653 = _T_189 | _T_652; // @[Lookup.scala 11:37]
  wire  _T_654 = _T_185 | _T_653; // @[Lookup.scala 11:37]
  wire  _T_655 = _T_181 | _T_654; // @[Lookup.scala 11:37]
  wire  _T_656 = _T_177 | _T_655; // @[Lookup.scala 11:37]
  wire  _T_657 = _T_173 | _T_656; // @[Lookup.scala 11:37]
  wire  _T_658 = _T_169 | _T_657; // @[Lookup.scala 11:37]
  wire  _T_659 = _T_165 | _T_658; // @[Lookup.scala 11:37]
  wire  _T_660 = _T_161 | _T_659; // @[Lookup.scala 11:37]
  wire  _T_661 = _T_157 | _T_660; // @[Lookup.scala 11:37]
  wire  _T_662 = _T_153 | _T_661; // @[Lookup.scala 11:37]
  wire  _T_663 = _T_149 | _T_662; // @[Lookup.scala 11:37]
  wire  _T_664 = _T_145 | _T_663; // @[Lookup.scala 11:37]
  wire  _T_665 = _T_141 | _T_664; // @[Lookup.scala 11:37]
  wire  _T_666 = _T_137 | _T_665; // @[Lookup.scala 11:37]
  wire  _T_667 = _T_133 | _T_666; // @[Lookup.scala 11:37]
  wire  _T_668 = _T_129 | _T_667; // @[Lookup.scala 11:37]
  wire  _T_669 = _T_125 | _T_668; // @[Lookup.scala 11:37]
  wire  _T_670 = _T_121 | _T_669; // @[Lookup.scala 11:37]
  wire  _T_671 = _T_117 ? 1'h0 : _T_670; // @[Lookup.scala 11:37]
  wire  _T_672 = _T_113 ? 1'h0 : _T_671; // @[Lookup.scala 11:37]
  wire  _T_673 = _T_109 ? 1'h0 : _T_672; // @[Lookup.scala 11:37]
  wire  _T_674 = _T_105 | _T_673; // @[Lookup.scala 11:37]
  wire  _T_675 = _T_101 | _T_674; // @[Lookup.scala 11:37]
  wire  _T_676 = _T_97 | _T_675; // @[Lookup.scala 11:37]
  wire  _T_677 = _T_93 | _T_676; // @[Lookup.scala 11:37]
  wire  cs0_2 = _T_89 | _T_677; // @[Lookup.scala 11:37]
  wire  _T_699 = _T_201 | _T_205; // @[Lookup.scala 11:37]
  wire  _T_700 = _T_197 | _T_699; // @[Lookup.scala 11:37]
  wire  _T_701 = _T_193 | _T_700; // @[Lookup.scala 11:37]
  wire  _T_702 = _T_189 | _T_701; // @[Lookup.scala 11:37]
  wire  _T_703 = _T_185 | _T_702; // @[Lookup.scala 11:37]
  wire  _T_704 = _T_181 | _T_703; // @[Lookup.scala 11:37]
  wire  _T_705 = _T_177 | _T_704; // @[Lookup.scala 11:37]
  wire  _T_706 = _T_173 | _T_705; // @[Lookup.scala 11:37]
  wire  _T_707 = _T_169 | _T_706; // @[Lookup.scala 11:37]
  wire  _T_708 = _T_165 | _T_707; // @[Lookup.scala 11:37]
  wire  _T_709 = _T_161 | _T_708; // @[Lookup.scala 11:37]
  wire  _T_710 = _T_157 | _T_709; // @[Lookup.scala 11:37]
  wire  _T_711 = _T_153 | _T_710; // @[Lookup.scala 11:37]
  wire  _T_712 = _T_149 | _T_711; // @[Lookup.scala 11:37]
  wire  _T_713 = _T_145 | _T_712; // @[Lookup.scala 11:37]
  wire  _T_714 = _T_141 | _T_713; // @[Lookup.scala 11:37]
  wire  _T_715 = _T_137 | _T_714; // @[Lookup.scala 11:37]
  wire  _T_716 = _T_133 | _T_715; // @[Lookup.scala 11:37]
  wire  _T_717 = _T_129 | _T_716; // @[Lookup.scala 11:37]
  wire  _T_718 = _T_125 | _T_717; // @[Lookup.scala 11:37]
  wire  _T_719 = _T_121 | _T_718; // @[Lookup.scala 11:37]
  wire  _T_720 = _T_117 ? 1'h0 : _T_719; // @[Lookup.scala 11:37]
  wire  _T_721 = _T_113 ? 1'h0 : _T_720; // @[Lookup.scala 11:37]
  wire  _T_722 = _T_109 ? 1'h0 : _T_721; // @[Lookup.scala 11:37]
  wire  _T_723 = _T_105 ? 1'h0 : _T_722; // @[Lookup.scala 11:37]
  wire  _T_724 = _T_101 ? 1'h0 : _T_723; // @[Lookup.scala 11:37]
  wire  _T_725 = _T_97 ? 1'h0 : _T_724; // @[Lookup.scala 11:37]
  wire  _T_726 = _T_93 ? 1'h0 : _T_725; // @[Lookup.scala 11:37]
  wire  _T_819 = _T_113 | _T_117; // @[Lookup.scala 11:37]
  wire  _T_820 = _T_109 | _T_819; // @[Lookup.scala 11:37]
  wire  _T_821 = _T_105 ? 1'h0 : _T_820; // @[Lookup.scala 11:37]
  wire  _T_822 = _T_101 ? 1'h0 : _T_821; // @[Lookup.scala 11:37]
  wire  _T_823 = _T_97 ? 1'h0 : _T_822; // @[Lookup.scala 11:37]
  wire  _T_824 = _T_93 ? 1'h0 : _T_823; // @[Lookup.scala 11:37]
  wire [2:0] _T_867 = _T_117 ? 3'h2 : 3'h0; // @[Lookup.scala 11:37]
  wire [2:0] _T_868 = _T_113 ? 3'h1 : _T_867; // @[Lookup.scala 11:37]
  wire [2:0] _T_869 = _T_109 ? 3'h3 : _T_868; // @[Lookup.scala 11:37]
  wire [2:0] _T_870 = _T_105 ? 3'h6 : _T_869; // @[Lookup.scala 11:37]
  wire [2:0] _T_871 = _T_101 ? 3'h2 : _T_870; // @[Lookup.scala 11:37]
  wire [2:0] _T_872 = _T_97 ? 3'h5 : _T_871; // @[Lookup.scala 11:37]
  wire [2:0] _T_873 = _T_93 ? 3'h1 : _T_872; // @[Lookup.scala 11:37]
  wire [2:0] _T_876 = _T_277 ? 3'h4 : 3'h0; // @[Lookup.scala 11:37]
  wire [2:0] _T_877 = _T_273 ? 3'h4 : _T_876; // @[Lookup.scala 11:37]
  wire [2:0] _T_878 = _T_269 ? 3'h4 : _T_877; // @[Lookup.scala 11:37]
  wire [2:0] _T_879 = _T_265 ? 3'h4 : _T_878; // @[Lookup.scala 11:37]
  wire [2:0] _T_880 = _T_261 ? 3'h4 : _T_879; // @[Lookup.scala 11:37]
  wire [2:0] _T_881 = _T_257 ? 3'h3 : _T_880; // @[Lookup.scala 11:37]
  wire [2:0] _T_882 = _T_253 ? 3'h3 : _T_881; // @[Lookup.scala 11:37]
  wire [2:0] _T_883 = _T_249 ? 3'h2 : _T_882; // @[Lookup.scala 11:37]
  wire [2:0] _T_884 = _T_245 ? 3'h1 : _T_883; // @[Lookup.scala 11:37]
  wire [2:0] _T_885 = _T_241 ? 3'h2 : _T_884; // @[Lookup.scala 11:37]
  wire [2:0] _T_886 = _T_237 ? 3'h1 : _T_885; // @[Lookup.scala 11:37]
  wire [2:0] _T_887 = _T_233 ? 3'h0 : _T_886; // @[Lookup.scala 11:37]
  wire [2:0] _T_888 = _T_229 ? 3'h0 : _T_887; // @[Lookup.scala 11:37]
  wire [2:0] _T_889 = _T_225 ? 3'h0 : _T_888; // @[Lookup.scala 11:37]
  wire [2:0] _T_890 = _T_221 ? 3'h0 : _T_889; // @[Lookup.scala 11:37]
  wire [2:0] _T_891 = _T_217 ? 3'h0 : _T_890; // @[Lookup.scala 11:37]
  wire [2:0] _T_892 = _T_213 ? 3'h0 : _T_891; // @[Lookup.scala 11:37]
  wire [2:0] _T_893 = _T_209 ? 3'h0 : _T_892; // @[Lookup.scala 11:37]
  wire [2:0] _T_894 = _T_205 ? 3'h0 : _T_893; // @[Lookup.scala 11:37]
  wire [2:0] _T_895 = _T_201 ? 3'h0 : _T_894; // @[Lookup.scala 11:37]
  wire [2:0] _T_896 = _T_197 ? 3'h0 : _T_895; // @[Lookup.scala 11:37]
  wire [2:0] _T_897 = _T_193 ? 3'h0 : _T_896; // @[Lookup.scala 11:37]
  wire [2:0] _T_898 = _T_189 ? 3'h0 : _T_897; // @[Lookup.scala 11:37]
  wire [2:0] _T_899 = _T_185 ? 3'h0 : _T_898; // @[Lookup.scala 11:37]
  wire [2:0] _T_900 = _T_181 ? 3'h0 : _T_899; // @[Lookup.scala 11:37]
  wire [2:0] _T_901 = _T_177 ? 3'h0 : _T_900; // @[Lookup.scala 11:37]
  wire [2:0] _T_902 = _T_173 ? 3'h0 : _T_901; // @[Lookup.scala 11:37]
  wire [2:0] _T_903 = _T_169 ? 3'h0 : _T_902; // @[Lookup.scala 11:37]
  wire [2:0] _T_904 = _T_165 ? 3'h0 : _T_903; // @[Lookup.scala 11:37]
  wire [2:0] _T_905 = _T_161 ? 3'h0 : _T_904; // @[Lookup.scala 11:37]
  wire [2:0] _T_906 = _T_157 ? 3'h0 : _T_905; // @[Lookup.scala 11:37]
  wire [2:0] _T_907 = _T_153 ? 3'h0 : _T_906; // @[Lookup.scala 11:37]
  wire [2:0] _T_908 = _T_149 ? 3'h0 : _T_907; // @[Lookup.scala 11:37]
  wire [2:0] _T_909 = _T_145 ? 3'h0 : _T_908; // @[Lookup.scala 11:37]
  wire [2:0] _T_910 = _T_141 ? 3'h0 : _T_909; // @[Lookup.scala 11:37]
  wire [2:0] _T_911 = _T_137 ? 3'h0 : _T_910; // @[Lookup.scala 11:37]
  wire [2:0] _T_912 = _T_133 ? 3'h0 : _T_911; // @[Lookup.scala 11:37]
  wire [2:0] _T_913 = _T_129 ? 3'h0 : _T_912; // @[Lookup.scala 11:37]
  wire [2:0] _T_914 = _T_125 ? 3'h0 : _T_913; // @[Lookup.scala 11:37]
  wire [2:0] _T_915 = _T_121 ? 3'h0 : _T_914; // @[Lookup.scala 11:37]
  wire [2:0] _T_916 = _T_117 ? 3'h0 : _T_915; // @[Lookup.scala 11:37]
  wire [2:0] _T_917 = _T_113 ? 3'h0 : _T_916; // @[Lookup.scala 11:37]
  wire [2:0] _T_918 = _T_109 ? 3'h0 : _T_917; // @[Lookup.scala 11:37]
  wire [2:0] _T_919 = _T_105 ? 3'h0 : _T_918; // @[Lookup.scala 11:37]
  wire [2:0] _T_920 = _T_101 ? 3'h0 : _T_919; // @[Lookup.scala 11:37]
  wire [2:0] _T_921 = _T_97 ? 3'h0 : _T_920; // @[Lookup.scala 11:37]
  wire [2:0] _T_922 = _T_93 ? 3'h0 : _T_921; // @[Lookup.scala 11:37]
  wire [2:0] cs0_7 = _T_89 ? 3'h0 : _T_922; // @[Lookup.scala 11:37]
  wire  _T_973 = cs_br_type == 4'h0; // @[cpath.scala 138:37]
  wire  _T_974 = cs_br_type == 4'h1; // @[cpath.scala 139:37]
  wire  _T_976 = ~io_dat_br_eq; // @[cpath.scala 139:54]
  wire [2:0] _T_977 = _T_976 ? 3'h1 : 3'h0; // @[cpath.scala 139:53]
  wire  _T_978 = cs_br_type == 4'h2; // @[cpath.scala 140:37]
  wire [2:0] _T_979 = io_dat_br_eq ? 3'h1 : 3'h0; // @[cpath.scala 140:53]
  wire  _T_980 = cs_br_type == 4'h3; // @[cpath.scala 141:37]
  wire  _T_982 = ~io_dat_br_lt; // @[cpath.scala 141:54]
  wire [2:0] _T_983 = _T_982 ? 3'h1 : 3'h0; // @[cpath.scala 141:53]
  wire  _T_984 = cs_br_type == 4'h4; // @[cpath.scala 142:37]
  wire  _T_986 = ~io_dat_br_ltu; // @[cpath.scala 142:54]
  wire [2:0] _T_987 = _T_986 ? 3'h1 : 3'h0; // @[cpath.scala 142:53]
  wire  _T_988 = cs_br_type == 4'h5; // @[cpath.scala 143:37]
  wire [2:0] _T_989 = io_dat_br_lt ? 3'h1 : 3'h0; // @[cpath.scala 143:53]
  wire  _T_990 = cs_br_type == 4'h6; // @[cpath.scala 144:37]
  wire [2:0] _T_991 = io_dat_br_ltu ? 3'h1 : 3'h0; // @[cpath.scala 144:53]
  wire  _T_992 = cs_br_type == 4'h7; // @[cpath.scala 145:37]
  wire  _T_993 = cs_br_type == 4'h8; // @[cpath.scala 146:37]
  wire [2:0] _T_994 = _T_993 ? 3'h3 : 3'h0; // @[cpath.scala 146:25]
  wire [2:0] _T_995 = _T_992 ? 3'h2 : _T_994; // @[cpath.scala 145:25]
  wire [2:0] _T_996 = _T_990 ? _T_991 : _T_995; // @[cpath.scala 144:25]
  wire [2:0] _T_997 = _T_988 ? _T_989 : _T_996; // @[cpath.scala 143:25]
  wire [2:0] _T_998 = _T_984 ? _T_987 : _T_997; // @[cpath.scala 142:25]
  wire [2:0] _T_999 = _T_980 ? _T_983 : _T_998; // @[cpath.scala 141:25]
  wire [2:0] _T_1000 = _T_978 ? _T_979 : _T_999; // @[cpath.scala 140:25]
  wire [2:0] _T_1001 = _T_974 ? _T_977 : _T_1000; // @[cpath.scala 139:25]
  wire [2:0] _T_1002 = _T_973 ? 3'h0 : _T_1001; // @[cpath.scala 138:25]
  reg  _T_1028; // @[cpath.scala 179:27]
  wire  take_evec = _T_1028 | io_dat_csr_eret; // @[cpath.scala 179:51]
  wire [2:0] ctrl_pc_sel = take_evec ? 3'h4 : _T_1002; // @[cpath.scala 137:25]
  wire  _T_1003 = ctrl_pc_sel == 3'h0; // @[cpath.scala 150:39]
  wire  _T_1005 = ~_T_1003; // @[cpath.scala 150:25]
  wire  _T_1009 = ~io_imem_resp_valid; // @[cpath.scala 159:29]
  wire [4:0] rs1_addr = io_imem_resp_bits_inst[19:15]; // @[cpath.scala 162:41]
  wire  _T_1014 = cs0_7 == 3'h2; // @[cpath.scala 163:30]
  wire  _T_1015 = cs0_7 == 3'h3; // @[cpath.scala 163:54]
  wire  _T_1016 = _T_1014 | _T_1015; // @[cpath.scala 163:40]
  wire  _T_1018 = rs1_addr == 5'h0; // @[cpath.scala 163:77]
  wire  csr_ren = _T_1016 & _T_1018; // @[cpath.scala 163:65]
  wire [2:0] csr_cmd = csr_ren ? 3'h5 : cs0_7; // @[cpath.scala 164:21]
  wire  _T_1025 = ~cs_inst_val; // @[cpath.scala 178:24]
  assign io_imem_req_valid = _T_1005 & io_imem_resp_valid; // @[cpath.scala 150:22]
  assign io_ctl_exe_kill = _T_1028 | io_dat_csr_eret; // @[cpath.scala 152:22]
  assign io_ctl_pc_sel = take_evec ? 3'h4 : _T_1002; // @[cpath.scala 153:22]
  assign io_ctl_brjmp_sel = _T_89 ? 1'h0 : _T_432; // @[cpath.scala 154:22]
  assign io_ctl_op1_sel = _T_89 ? 2'h0 : _T_481; // @[cpath.scala 155:22]
  assign io_ctl_op2_sel = _T_89 ? 2'h1 : _T_530; // @[cpath.scala 156:22]
  assign io_ctl_alu_fun = _T_89 ? 4'h0 : _T_579; // @[cpath.scala 157:22]
  assign io_ctl_wb_sel = _T_89 ? 2'h1 : _T_628; // @[cpath.scala 158:22]
  assign io_ctl_rf_wen = _T_1009 ? 1'h0 : cs0_2; // @[cpath.scala 159:22]
  assign io_ctl_bypassable = _T_89 ? 1'h0 : _T_726; // @[cpath.scala 160:22]
  assign io_ctl_csr_cmd = _T_1009 ? 3'h0 : csr_cmd; // @[cpath.scala 165:22]
  assign io_ctl_dmem_fcn = _T_89 ? 1'h0 : _T_824; // @[cpath.scala 172:22]
  assign io_ctl_dmem_typ = _T_89 ? 3'h3 : _T_873; // @[cpath.scala 173:22]
  assign io_ctl_exception = _T_1025 & io_imem_resp_valid; // @[cpath.scala 178:21]
  assign _GEN_92_0 = 32'h3013 == _T_88;
  assign _GEN_52_0 = 32'h4013 == _T_88;
  assign _GEN_305_0 = cs_br_type == 4'h5;
  assign _GEN_200_0 = 32'h40000033 == _T_164;
  assign _GEN_149_0 = 32'h67 == _T_88;
  assign _GEN_25_0 = 32'h7013 == _T_88;
  assign _GEN_248_0 = 32'h10500073 == io_imem_resp_bits_inst;
  assign _GEN_107_0 = 32'h67 == _T_88;
  assign _GEN_134_0 = 32'h1003 == _T_88;
  assign _GEN_206_0 = 32'h3013 == _T_88;
  assign _GEN_40_0 = 32'h6033 == _T_164;
  assign _GEN_233_0 = 32'h5003 == _T_88;
  assign _GEN_128_0 = 32'h37 == _T_120;
  assign _GEN_191_0 = 32'h67 == _T_88;
  assign _GEN_227_0 = 32'h1023 == _T_88;
  assign _GEN_113_0 = 32'h7033 == _T_164;
  assign _GEN_46_0 = 32'h1033 == _T_164;
  assign _GEN_299_0 = ~io_dat_br_ltu;
  assign _GEN_73_0 = 32'h7063 == _T_88;
  assign _GEN_212_0 = 32'h37 == _T_120;
  assign _GEN_31_0 = 32'h2023 == _T_88;
  assign _GEN_311_0 = _T_1028 | io_dat_csr_eret;
  assign _GEN_67_0 = 32'h2073 == _T_88;
  assign _GEN_320_0 = 32'h2003 == _T_88;
  assign _GEN_215_0 = 32'h23 == _T_88;
  assign _GEN_221_0 = 32'h6063 == _T_88;
  assign _GEN_101_0 = 32'h23 == _T_88;
  assign _GEN_110_0 = 32'h40005033 == _T_164;
  assign _GEN_283_0 = 32'h6013 == _T_88;
  assign _GEN_314_0 = 32'h2003 == _T_88;
  assign _GEN_178_0 = 32'h3 == _T_88;
  assign _GEN_209_0 = 32'h6013 == _T_88;
  assign _GEN_28_0 = 32'h17 == _T_120;
  assign _GEN_277_0 = 32'h5013 == _T_152;
  assign _GEN_55_0 = 32'h13 == _T_88;
  assign _GEN_194_0 = 32'h40005033 == _T_164;
  assign _GEN_13_0 = 32'h3033 == _T_164;
  assign _GEN_49_0 = 32'h1013 == _T_152;
  assign _GEN_116_0 = 32'h40000033 == _T_164;
  assign _GEN_7_0 = 32'h6f == _T_120;
  assign _GEN_34_0 = 32'h4003 == _T_88;
  assign _GEN_122_0 = 32'h3013 == _T_88;
  assign _GEN_308_0 = cs_br_type == 4'h2;
  assign _GEN_95_0 = 32'h6013 == _T_88;
  assign _GEN_230_0 = 32'h1023 == _T_88;
  assign _GEN_293_0 = 32'h4003 == _T_88;
  assign _GEN_184_0 = 32'h5073 == _T_88;
  assign _GEN_1_2 = 32'h4063 == _T_88;
  assign _GEN_197_0 = 32'h7033 == _T_164;
  assign _GEN_187_0 = 32'h7063 == _T_88;
  assign _GEN_104_0 = 32'h1003 == _T_88;
  assign _GEN_265_0 = 32'h67 == _T_88;
  assign _GEN_296_0 = ~io_dat_br_eq;
  assign _GEN_160_0 = 32'h1033 == _T_164;
  assign _GEN_172_0 = 32'h1023 == _T_88;
  assign _GEN_203_0 = 32'h5013 == _T_152;
  assign _GEN_271_0 = 32'h7033 == _T_164;
  assign _GEN_37_0 = 32'h5033 == _T_164;
  assign _GEN_166_0 = 32'h4013 == _T_88;
  assign _GEN_280_0 = 32'h3013 == _T_88;
  assign _GEN_286_0 = 32'h37 == _T_120;
  assign _GEN_22_1 = 32'h2013 == _T_88;
  assign _GEN_302_0 = cs_br_type == 4'h8;
  assign _GEN_16_2 = 32'h33 == _T_164;
  assign _GEN_10_2 = 32'h4033 == _T_164;
  assign _GEN_259_0 = 32'h6063 == _T_88;
  assign _GEN_98_0 = 32'h37 == _T_120;
  assign _GEN_19_1 = 32'h40005013 == _T_152;
  assign _GEN_148_0 = 32'h63 == _T_88;
  assign _GEN_87_0 = 32'h33 == _T_164;
  assign _GEN_274_0 = 32'h40000033 == _T_164;
  assign _GEN_232_0 = 32'h2023 == _T_88;
  assign _GEN_190_0 = 32'h63 == _T_88;
  assign _GEN_154_0 = 32'h6033 == _T_164;
  assign _GEN_289_0 = 32'h23 == _T_88;
  assign _GEN_181_0 = 32'h2073 == _T_88;
  assign _GEN_253_0 = 32'h7073 == _T_88;
  assign _GEN_72_0 = 32'h4063 == _T_88;
  assign _GEN_175_0 = 32'h5003 == _T_88;
  assign _GEN_169_0 = 32'h13 == _T_88;
  assign _GEN_4_1 = 32'h1063 == _T_88;
  assign _GEN_247_0 = 32'h3 == _T_88;
  assign _GEN_268_0 = 32'h40005033 == _T_164;
  assign _GEN_214_0 = 32'h1023 == _T_88;
  assign _GEN_250_0 = 32'h7b200073 == io_imem_resp_bits_inst;
  assign _GEN_241_0 = 32'h1023 == _T_88;
  assign _GEN_142_0 = 32'h5073 == _T_88;
  assign _GEN_136_0 = 32'h3 == _T_88;
  assign _GEN_235_0 = 32'h4003 == _T_88;
  assign _GEN_262_0 = 32'h5063 == _T_88;
  assign _GEN_54_0 = 32'h7013 == _T_88;
  assign _GEN_313_0 = _T_1028 | io_dat_csr_eret;
  assign _GEN_69_0 = 32'h6073 == _T_88;
  assign _GEN_157_0 = 32'h2033 == _T_164;
  assign _GEN_75_0 = 32'h1063 == _T_88;
  assign _GEN_90_0 = 32'h40005013 == _T_152;
  assign _GEN_163_0 = 32'h1013 == _T_152;
  assign _GEN_130_0 = 32'h1023 == _T_88;
  assign _GEN_229_0 = 32'h2023 == _T_88;
  assign _GEN_121_0 = 32'h1013 == _T_152;
  assign _GEN_256_0 = 32'h1073 == _T_88;
  assign _GEN_81_0 = 32'h4033 == _T_164;
  assign _GEN_57_0 = 32'h17 == _T_120;
  assign _GEN_145_0 = 32'h7063 == _T_88;
  assign _GEN_223_0 = 32'h7063 == _T_88;
  assign _GEN_118_0 = 32'h1033 == _T_164;
  assign _GEN_322_0 = 32'h2003 == _T_88;
  assign _GEN_244_0 = 32'h5003 == _T_88;
  assign _GEN_124_0 = 32'h4013 == _T_88;
  assign _GEN_103_0 = 32'h5003 == _T_88;
  assign _GEN_238_0 = 32'h1003 == _T_88;
  assign _GEN_63_0 = 32'h4003 == _T_88;
  assign _GEN_151_0 = 32'h5033 == _T_164;
  assign _GEN_202_0 = 32'h1033 == _T_164;
  assign _GEN_196_0 = 32'h6033 == _T_164;
  assign _GEN_295_0 = 32'h2003 == _T_88;
  assign _GEN_301_0 = io_dat_br_ltu;
  assign _GEN_310_0 = cs_br_type == 4'h0;
  assign _GEN_78_0 = 32'h6f == _T_120;
  assign _GEN_84_0 = 32'h3033 == _T_164;
  assign _GEN_217_0 = 32'h5003 == _T_88;
  assign _GEN_36_0 = 32'h2003 == _T_88;
  assign _GEN_42_0 = 32'h3033 == _T_164;
  assign _GEN_316_0 = 32'h2003 == _T_88;
  assign _GEN_139_0 = 32'h2073 == _T_88;
  assign _GEN_18_1 = 32'h5013 == _T_152;
  assign _GEN_226_0 = 32'h63 == _T_88;
  assign _GEN_106_0 = 32'h3 == _T_88;
  assign _GEN_51_0 = 32'h2013 == _T_88;
  assign _GEN_45_0 = 32'h33 == _T_164;
  assign _GEN_319_0 = ~io_imem_resp_valid;
  assign _GEN_39_0 = 32'h4033 == _T_164;
  assign _GEN_66_0 = 32'h3073 == _T_88;
  assign _GEN_24_0 = 32'h6013 == _T_88;
  assign _GEN_112_0 = 32'h6033 == _T_164;
  assign _GEN_211_0 = 32'h13 == _T_88;
  assign _GEN_220_0 = 32'h3 == _T_88;
  assign _GEN_133_0 = 32'h5003 == _T_88;
  assign _GEN_127_0 = 32'h13 == _T_88;
  assign _GEN_288_1 = 32'h1023 == _T_88;
  assign _GEN_91_0 = 32'h1013 == _T_152;
  assign _GEN_205_0 = 32'h1013 == _T_152;
  assign _GEN_100_0 = 32'h1023 == _T_88;
  assign _GEN_304_0 = cs_br_type == 4'h6;
  assign _GEN_60_0 = 32'h2023 == _T_88;
  assign _GEN_298_0 = ~io_dat_br_lt;
  assign _GEN_189_0 = 32'h1063 == _T_88;
  assign _GEN_199_0 = 32'h2033 == _T_164;
  assign _GEN_177_0 = 32'h4003 == _T_88;
  assign _GEN_12_2 = 32'h7033 == _T_164;
  assign _GEN_94_0 = 32'h4013 == _T_88;
  assign _GEN_162_0 = 32'h40005013 == _T_152;
  assign _GEN_193_0 = 32'h5033 == _T_164;
  assign _GEN_208_0 = 32'h4013 == _T_88;
  assign _GEN_261_0 = 32'h7063 == _T_88;
  assign _GEN_115_0 = 32'h2033 == _T_164;
  assign _GEN_27_0 = 32'h37 == _T_120;
  assign _GEN_270_0 = 32'h6033 == _T_164;
  assign _GEN_183_0 = 32'h6073 == _T_88;
  assign _GEN_33_0 = 32'h1003 == _T_88;
  assign _GEN_276_0 = 32'h1033 == _T_164;
  assign _GEN_282_1 = 32'h4013 == _T_88;
  assign _GEN_292_0 = 32'h1003 == _T_88;
  assign _GEN_48_0 = 32'h40005013 == _T_152;
  assign _GEN_6_2 = 32'h67 == _T_88;
  assign _GEN_307_0 = cs_br_type == 4'h3;
  assign _GEN_109_0 = 32'h5033 == _T_164;
  assign _GEN_21_1 = 32'h3013 == _T_88;
  assign _GEN_15_3 = 32'h40000033 == _T_164;
  assign _GEN_30_0 = 32'h23 == _T_88;
  assign _GEN_83_0 = 32'h7033 == _T_164;
  assign _GEN_171_0 = 32'h17 == _T_120;
  assign _GEN_186_0 = 32'h4063 == _T_88;
  assign _GEN_144_0 = 32'h4063 == _T_88;
  assign _GEN_279_1 = 32'h1013 == _T_152;
  assign _GEN_97_0 = 32'h13 == _T_88;
  assign _GEN_264_0 = 32'h63 == _T_88;
  assign _GEN_165_0 = 32'h2013 == _T_88;
  assign _GEN_159_0 = 32'h33 == _T_164;
  assign _GEN_258_0 = 32'h5073 == _T_88;
  assign _GEN_285_1 = 32'h13 == _T_88;
  assign _GEN_180_0 = 32'h3073 == _T_88;
  assign _GEN_9_3 = 32'h40005033 == _T_164;
  assign _GEN_243_0 = 32'h2023 == _T_88;
  assign _GEN_77_0 = 32'h67 == _T_88;
  assign _GEN_174_0 = 32'h2023 == _T_88;
  assign _GEN_225_0 = 32'h1063 == _T_88;
  assign _GEN_252_0 = 32'h73 == io_imem_resp_bits_inst;
  assign _GEN_132_0 = 32'h2023 == _T_88;
  assign _GEN_147_1 = 32'h1063 == _T_88;
  assign _GEN_240_0 = 32'h3 == _T_88;
  assign _GEN_65_0 = 32'h7073 == _T_88;
  assign _GEN_273_0 = 32'h2033 == _T_164;
  assign _GEN_59_0 = 32'h23 == _T_88;
  assign _GEN_231_0 = 32'h23 == _T_88;
  assign _GEN_86_0 = 32'h40000033 == _T_164;
  assign _GEN_80_0 = 32'h40005033 == _T_164;
  assign _GEN_3_2 = 32'h5063 == _T_88;
  assign _GEN_246_0 = 32'h4003 == _T_88;
  assign _GEN_71_0 = 32'h6063 == _T_88;
  assign _GEN_153_0 = 32'h4033 == _T_164;
  assign _GEN_168_0 = 32'h7013 == _T_88;
  assign _GEN_267_0 = 32'h5033 == _T_164;
  assign _GEN_126_0 = 32'h7013 == _T_88;
  assign _GEN_213_0 = 32'h17 == _T_120;
  assign _GEN_255_0 = 32'h2073 == _T_88;
  assign _GEN_156_0 = 32'h3033 == _T_164;
  assign _GEN_150_0 = 32'h6f == _T_120;
  assign _GEN_114_0 = 32'h3033 == _T_164;
  assign _GEN_228_0 = 32'h23 == _T_88;
  assign _GEN_141_0 = 32'h6073 == _T_88;
  assign _GEN_108_0 = 32'h6f == _T_120;
  assign _GEN_249_0 = 32'h100073 == io_imem_resp_bits_inst;
  assign _GEN_312_1 = _T_1016 & _T_1018;
  assign _GEN_68_0 = 32'h1073 == _T_88;
  assign _GEN_74_0 = 32'h5063 == _T_88;
  assign _GEN_207_0 = 32'h2013 == _T_88;
  assign _GEN_234_0 = 32'h1003 == _T_88;
  assign _GEN_306_1 = cs_br_type == 4'h4;
  assign _GEN_129_0 = 32'h17 == _T_120;
  assign _GEN_89_0 = 32'h5013 == _T_152;
  assign _GEN_47_0 = 32'h5013 == _T_152;
  assign _GEN_53_0 = 32'h6013 == _T_88;
  assign _GEN_135_0 = 32'h4003 == _T_88;
  assign _GEN_222_0 = 32'h4063 == _T_88;
  assign _GEN_29_0 = 32'h1023 == _T_88;
  assign _GEN_41_0 = 32'h7033 == _T_164;
  assign _GEN_56_0 = 32'h37 == _T_120;
  assign _GEN_195_0 = 32'h4033 == _T_164;
  assign _GEN_237_0 = 32'h5003 == _T_88;
  assign _GEN_102_0 = 32'h2023 == _T_88;
  assign _GEN_62_0 = 32'h1003 == _T_88;
  assign _GEN_35_0 = 32'h3 == _T_88;
  assign _GEN_123_0 = 32'h2013 == _T_88;
  assign _GEN_117_0 = 32'h33 == _T_164;
  assign _GEN_321_0 = ~io_imem_resp_valid;
  assign _GEN_216_0 = 32'h2023 == _T_88;
  assign _GEN_294_1 = 32'h3 == _T_88;
  assign _GEN_50_0 = 32'h3013 == _T_88;
  assign _GEN_138_0 = 32'h3073 == _T_88;
  assign _GEN_201_0 = 32'h33 == _T_164;
  assign _GEN_210_0 = 32'h7013 == _T_88;
  assign _GEN_96_0 = 32'h7013 == _T_88;
  assign _GEN_315_0 = 32'h2003 == _T_88;
  assign _GEN_309_0 = cs_br_type == 4'h1;
  assign _GEN_17_1 = 32'h1033 == _T_164;
  assign _GEN_105_0 = 32'h4003 == _T_88;
  assign _GEN_303_0 = cs_br_type == 4'h7;
  assign _GEN_204_0 = 32'h40005013 == _T_152;
  assign _GEN_318_1 = 32'h2003 == _T_88;
  assign _GEN_173_0 = 32'h23 == _T_88;
  assign _GEN_198_0 = 32'h3033 == _T_164;
  assign _GEN_23_1 = 32'h4013 == _T_88;
  assign _GEN_272_1 = 32'h3033 == _T_164;
  assign _GEN_120_0 = 32'h40005013 == _T_152;
  assign _GEN_188_0 = 32'h5063 == _T_88;
  assign _GEN_44_0 = 32'h40000033 == _T_164;
  assign _GEN_287_1 = 32'h17 == _T_120;
  assign _GEN_297_0 = io_dat_br_eq;
  assign _GEN_2_2 = 32'h7063 == _T_88;
  assign _GEN_99_0 = 32'h17 == _T_120;
  assign _GEN_38_0 = 32'h40005033 == _T_164;
  assign _GEN_111_0 = 32'h4033 == _T_164;
  assign _GEN_219_0 = 32'h4003 == _T_88;
  assign _GEN_26_0 = 32'h13 == _T_88;
  assign _GEN_176_0 = 32'h1003 == _T_88;
  assign _GEN_182_0 = 32'h1073 == _T_88;
  assign _GEN_290_1 = 32'h2023 == _T_88;
  assign _GEN_0_2 = 32'h6063 == _T_88;
  assign _GEN_32_0 = 32'h5003 == _T_88;
  assign _GEN_161_0 = 32'h5013 == _T_152;
  assign _GEN_275_1 = 32'h33 == _T_164;
  assign _GEN_170_0 = 32'h37 == _T_120;
  assign _GEN_192_0 = 32'h6f == _T_120;
  assign _GEN_20_1 = 32'h1013 == _T_152;
  assign _GEN_269_1 = 32'h4033 == _T_164;
  assign _GEN_281_1 = 32'h2013 == _T_88;
  assign _GEN_291_1 = 32'h5003 == _T_88;
  assign _GEN_155_0 = 32'h7033 == _T_164;
  assign _GEN_88_0 = 32'h1033 == _T_164;
  assign _GEN_300_1 = io_dat_br_lt;
  assign _GEN_11_3 = 32'h6033 == _T_164;
  assign _GEN_5_3 = 32'h63 == _T_88;
  assign _GEN_254_1 = 32'h3073 == _T_88;
  assign _GEN_93_0 = 32'h2013 == _T_88;
  assign _GEN_14_2 = 32'h2033 == _T_164;
  assign _GEN_257_1 = 32'h6073 == _T_88;
  assign _GEN_82_0 = 32'h6033 == _T_164;
  assign _GEN_8_2 = 32'h5033 == _T_164;
  assign _GEN_278_1 = 32'h40005013 == _T_152;
  assign _GEN_70_0 = 32'h5073 == _T_88;
  assign _GEN_158_0 = 32'h40000033 == _T_164;
  assign _GEN_236_1 = 32'h3 == _T_88;
  assign _GEN_185_0 = 32'h6063 == _T_88;
  assign _GEN_61_0 = 32'h5003 == _T_88;
  assign _GEN_143_0 = 32'h6063 == _T_88;
  assign _GEN_284_1 = 32'h7013 == _T_88;
  assign _GEN_179_0 = 32'h7073 == _T_88;
  assign _GEN_242_1 = 32'h23 == _T_88;
  assign _GEN_137_0 = 32'h7073 == _T_88;
  assign _GEN_76_0 = 32'h63 == _T_88;
  assign _GEN_164_0 = 32'h3013 == _T_88;
  assign _GEN_263_1 = 32'h1063 == _T_88;
  assign _GEN_167_0 = 32'h6013 == _T_88;
  assign _GEN_43_0 = 32'h2033 == _T_164;
  assign _GEN_266_1 = 32'h6f == _T_120;
  assign _GEN_131_0 = 32'h23 == _T_88;
  assign _GEN_125_0 = 32'h6013 == _T_88;
  assign _GEN_317_1 = 32'h2003 == _T_88;
  assign _GEN_224_0 = 32'h5063 == _T_88;
  assign _GEN_119_0 = 32'h5013 == _T_152;
  assign _GEN_239_1 = 32'h4003 == _T_88;
  assign _GEN_152_1 = 32'h40005033 == _T_164;
  assign _GEN_146_1 = 32'h5063 == _T_88;
  assign _GEN_245_1 = 32'h1003 == _T_88;
  assign _GEN_323_1 = 32'h2003 == _T_88;
  assign _GEN_79_0 = 32'h5033 == _T_164;
  assign _GEN_218_0 = 32'h1003 == _T_88;
  assign _GEN_64_0 = 32'h3 == _T_88;
  assign _GEN_58_0 = 32'h1023 == _T_88;
  assign _GEN_251_1 = 32'h30200073 == io_imem_resp_bits_inst;
  assign _GEN_260_1 = 32'h4063 == _T_88;
  assign _GEN_140_0 = 32'h1073 == _T_88;
  assign _GEN_85_0 = 32'h2033 == _T_164;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1028 = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      _T_1028 <= 1'h0;
    end else begin
      _T_1028 <= io_ctl_exception;
    end
  end
endmodule
module ALU(
  input  [3:0]  io_fn,
  input  [31:0] io_in2,
  input  [31:0] io_in1,
  output [31:0] io_out,
  output [31:0] io_adder_out,
  output        _GEN_16_0,
  output        _GEN_10_0,
  output        _GEN_15_1,
  output        _GEN_18_0,
  output        _GEN_12_1,
  output        _GEN_9_1,
  output        _GEN_8_1,
  output        _GEN_11_2,
  output        _GEN_17_0,
  output        _GEN_14_0,
  output        _GEN_13_3
);
  wire [31:0] _T_13 = 32'h0 - io_in2; // @[alu.scala 50:40]
  wire [31:0] _T_14 = io_fn[3] ? _T_13 : io_in2; // @[alu.scala 50:25]
  wire [31:0] sum = io_in1 + _T_14; // @[alu.scala 50:20]
  wire  _T_18 = io_in1[31] == io_in2[31]; // @[alu.scala 53:32]
  wire  _T_23 = io_fn[1] ? io_in2[31] : io_in1[31]; // @[alu.scala 54:18]
  wire  less = _T_18 ? sum[31] : _T_23; // @[alu.scala 53:19]
  wire [4:0] shamt = io_in2[4:0]; // @[alu.scala 58:21]
  wire  _T_24 = io_fn == 4'h5; // @[alu.scala 60:24]
  wire  _T_25 = io_fn == 4'hb; // @[alu.scala 60:46]
  wire  _T_26 = _T_24 | _T_25; // @[alu.scala 60:37]
  wire [31:0] _T_32 = {{16'd0}, io_in1[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_34 = {io_in1[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_36 = _T_34 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_37 = _T_32 | _T_36; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_0 = {{8'd0}, _T_37[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_42 = _GEN_0 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_44 = {_T_37[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_46 = _T_44 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_47 = _T_42 | _T_46; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1 = {{4'd0}, _T_47[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_52 = _GEN_1 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_54 = {_T_47[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_56 = _T_54 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_57 = _T_52 | _T_56; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_2 = {{2'd0}, _T_57[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_62 = _GEN_2 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_64 = {_T_57[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_66 = _T_64 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_67 = _T_62 | _T_66; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_3 = {{1'd0}, _T_67[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_72 = _GEN_3 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_74 = {_T_67[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_76 = _T_74 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] _T_77 = _T_72 | _T_76; // @[Bitwise.scala 103:39]
  wire [31:0] shin = _T_26 ? io_in1 : _T_77; // @[alu.scala 60:17]
  wire  _T_80 = io_fn[3] & shin[31]; // @[alu.scala 61:35]
  wire [32:0] _T_82 = {_T_80,shin};
  wire [32:0] _T_83 = $signed(_T_82) >>> shamt; // @[alu.scala 61:61]
  wire [31:0] shout_r = _T_83[31:0]; // @[alu.scala 61:70]
  wire [31:0] _T_89 = {{16'd0}, shout_r[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_91 = {shout_r[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_93 = _T_91 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_94 = _T_89 | _T_93; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_4 = {{8'd0}, _T_94[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_99 = _GEN_4 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_101 = {_T_94[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_103 = _T_101 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_104 = _T_99 | _T_103; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_5 = {{4'd0}, _T_104[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_109 = _GEN_5 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_111 = {_T_104[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_113 = _T_111 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_114 = _T_109 | _T_113; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_6 = {{2'd0}, _T_114[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_119 = _GEN_6 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_121 = {_T_114[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_123 = _T_121 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_124 = _T_119 | _T_123; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_7 = {{1'd0}, _T_124[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_129 = _GEN_7 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_131 = {_T_124[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_133 = _T_131 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] shout_l = _T_129 | _T_133; // @[Bitwise.scala 103:39]
  wire  _T_134 = io_fn == 4'h7; // @[alu.scala 65:15]
  wire [31:0] _T_135 = io_in1 & io_in2; // @[alu.scala 65:35]
  wire  _T_136 = io_fn == 4'h6; // @[alu.scala 66:15]
  wire [31:0] _T_137 = io_in1 | io_in2; // @[alu.scala 66:35]
  wire  _T_138 = io_fn == 4'h4; // @[alu.scala 67:15]
  wire [31:0] _T_139 = io_in1 ^ io_in2; // @[alu.scala 67:35]
  wire [31:0] _T_140 = _T_138 ? _T_139 : io_in1; // @[alu.scala 67:8]
  wire [31:0] _T_141 = _T_136 ? _T_137 : _T_140; // @[alu.scala 66:8]
  wire [31:0] bitwise_logic = _T_134 ? _T_135 : _T_141; // @[alu.scala 65:8]
  wire  _T_142 = io_fn == 4'h0; // @[alu.scala 71:15]
  wire  _T_143 = io_fn == 4'ha; // @[alu.scala 71:36]
  wire  _T_144 = _T_142 | _T_143; // @[alu.scala 71:27]
  wire  _T_145 = io_fn == 4'hc; // @[alu.scala 72:15]
  wire  _T_146 = io_fn == 4'he; // @[alu.scala 72:36]
  wire  _T_147 = _T_145 | _T_146; // @[alu.scala 72:27]
  wire  _T_151 = io_fn == 4'h1; // @[alu.scala 74:15]
  wire [31:0] _T_152 = _T_151 ? shout_l : bitwise_logic; // @[alu.scala 74:8]
  wire [31:0] _T_153 = _T_26 ? shout_r : _T_152; // @[alu.scala 73:8]
  wire [31:0] _T_154 = _T_147 ? {{31'd0}, less} : _T_153; // @[alu.scala 72:8]
  assign io_out = _T_144 ? sum : _T_154; // @[alu.scala 77:10]
  assign io_adder_out = io_in1 + _T_14; // @[alu.scala 78:16]
  assign _GEN_16_0 = _T_24 | _T_25;
  assign _GEN_10_0 = io_in1[31] == io_in2[31];
  assign _GEN_15_1 = io_fn == 4'h1;
  assign _GEN_18_0 = _T_142 | _T_143;
  assign _GEN_12_1 = io_fn == 4'h4;
  assign _GEN_9_1 = io_fn[1];
  assign _GEN_8_1 = io_fn[3];
  assign _GEN_11_2 = _T_24 | _T_25;
  assign _GEN_17_0 = _T_145 | _T_146;
  assign _GEN_14_0 = io_fn == 4'h7;
  assign _GEN_13_3 = io_fn == 4'h6;
endmodule
module CSRFile(
  input         metaReset,
  input         clock,
  input         reset,
  input  [2:0]  io_rw_cmd,
  output [31:0] io_rw_rdata,
  input  [31:0] io_rw_wdata,
  output        io_eret,
  input  [11:0] io_decode_csr,
  output        io_status_debug,
  output [1:0]  io_status_prv,
  output        io_status_sd,
  output [7:0]  io_status_zero1,
  output        io_status_tsr,
  output        io_status_tw,
  output        io_status_tvm,
  output        io_status_mxr,
  output        io_status_sum,
  output        io_status_mprv,
  output [1:0]  io_status_xs,
  output [1:0]  io_status_fs,
  output [1:0]  io_status_mpp,
  output [1:0]  io_status_hpp,
  output        io_status_spp,
  output        io_status_mpie,
  output        io_status_hpie,
  output        io_status_spie,
  output        io_status_upie,
  output        io_status_mie,
  output        io_status_hie,
  output        io_status_sie,
  output        io_status_uie,
  output [31:0] io_evec,
  input         io_exception,
  input         io_retire,
  input  [31:0] io_pc,
  output        _GEN_411_0,
  output        _GEN_405_0,
  output        _GEN_426_0,
  output        _GEN_291_0,
  output        _GEN_306_0,
  output        _GEN_384_0,
  output        _GEN_327_0,
  output        _GEN_390_0,
  output        _GEN_285_0,
  output        _GEN_318_0,
  output        _GEN_312_0,
  output        _GEN_399_0,
  output        _GEN_387_0,
  output        _GEN_300_0,
  output        _GEN_279_0,
  output        _GEN_269_0,
  output        _GEN_378_0,
  output        _GEN_368_0,
  output        _GEN_377_0,
  output        _GEN_294_0,
  output        _GEN_393_0,
  output        _GEN_362_0,
  output        _GEN_461_0,
  output        _GEN_263_0,
  output        _GEN_449_0,
  output        _GEN_288_0,
  output        _GEN_245_0,
  output        _GEN_272_0,
  output        _GEN_381_0,
  output        _GEN_371_0,
  output        _GEN_266_0,
  output        _GEN_344_0,
  output        _GEN_282_0,
  output        _GEN_443_0,
  output        _GEN_251_0,
  output        _GEN_350_0,
  output        _GEN_365_0,
  output        _GEN_15_0,
  output        _GEN_152_0,
  output        _GEN_446_0,
  output        _GEN_332_0,
  output        _GEN_326_0,
  output        _GEN_359_0,
  output        _GEN_458_0,
  output        _GEN_452_0,
  output        _GEN_347_0,
  output        _GEN_425_0,
  output        _GEN_239_0,
  output        _GEN_431_0,
  output        _GEN_254_0,
  output        _GEN_353_0,
  output        _GEN_260_0,
  output        _GEN_275_0,
  output        _GEN_338_0,
  output        _GEN_374_0,
  output        _GEN_242_0,
  output        _GEN_455_0,
  output        _GEN_413_0,
  output        _GEN_236_0,
  output        _GEN_335_0,
  output        _GEN_434_0,
  output        _GEN_248_1,
  output        _GEN_257_0,
  output        _GEN_320_1,
  output        _GEN_356_0,
  output        _GEN_419_0,
  output        _GEN_314_1,
  output        _GEN_341_0,
  output        _GEN_440_0,
  output        _GEN_299_1,
  output        _GEN_398_0,
  output        _GEN_407_0,
  output        _GEN_149_1,
  output        _GEN_416_0,
  output        _GEN_281_0,
  output        _GEN_380_0,
  output        _GEN_296_1,
  output        _GEN_422_0,
  output        _GEN_329_0,
  output        _GEN_6_1,
  output        _GEN_437_0,
  output        _GEN_302_1,
  output        _GEN_401_0,
  output        _GEN_395_0,
  output        _GEN_428_0,
  output        _GEN_308_1,
  output        _GEN_323_0,
  output        _GEN_317_0,
  output        _GEN_404_0,
  output        _GEN_290_0,
  output        _GEN_367_0,
  output        _GEN_284_0,
  output        _GEN_274_1,
  output        _GEN_383_0,
  output        _GEN_373_0,
  output        _GEN_410_0,
  output        _GEN_305_1,
  output        _GEN_311_1,
  output        _GEN_389_0,
  output        _GEN_268_1,
  output        _GEN_376_0,
  output        _GEN_454_0,
  output        _GEN_293_1,
  output        _GEN_392_0,
  output        _GEN_361_0,
  output        _GEN_287_0,
  output        _GEN_256_1,
  output        _GEN_460_0,
  output        _GEN_278_0,
  output        _GEN_355_0,
  output        _GEN_386_0,
  output        _GEN_277_1,
  output        _GEN_262_1,
  output        _GEN_244_1,
  output        _GEN_448_0,
  output        _GEN_442_0,
  output        _GEN_457_0,
  output        _GEN_337_0,
  output        _GEN_364_0,
  output        _GEN_328_0,
  output        _GEN_463_0,
  output        _GEN_436_0,
  output        _GEN_370_0,
  output        _GEN_250_1,
  output        _GEN_265_1,
  output        _GEN_271_1,
  output        _GEN_349_0,
  output        _GEN_343_0,
  output        _GEN_147_0,
  output        _GEN_352_0,
  output        _GEN_247_1,
  output        _GEN_325_0,
  output        _GEN_151_1,
  output        _GEN_238_1,
  output        _GEN_451_0,
  output        _GEN_346_0,
  output        _GEN_409_0,
  output        _GEN_253_1,
  output        _GEN_331_0,
  output        _GEN_11_1,
  output        _GEN_430_0,
  output        _GEN_424_0,
  output        _GEN_445_0,
  output        _GEN_310_1,
  output        _GEN_259_1,
  output        _GEN_358_0,
  output        _GEN_334_0,
  output        _GEN_412_0,
  output        _GEN_418_0,
  output        _GEN_427_0,
  output        _GEN_313_1,
  output        _GEN_292_1,
  output        _GEN_241_1,
  output        _GEN_340_0,
  output        _GEN_235_1,
  output        _GEN_439_0,
  output        _GEN_298_1,
  output        _GEN_307_1,
  output        _GEN_406_0,
  output        _GEN_433_0,
  output        _GEN_319_1,
  output        _GEN_391_0,
  output        _GEN_400_0,
  output        _GEN_415_0,
  output        _GEN_295_1,
  output        _GEN_270_1,
  output        _GEN_322_1,
  output        _GEN_421_0,
  output        _GEN_280_1,
  output        _GEN_379_0,
  output        _GEN_394_0,
  output        _GEN_369_0,
  output        _GEN_5_2,
  output        _GEN_316_1,
  output        _GEN_301_1,
  output        _GEN_283_1,
  output        _GEN_273_1,
  output        _GEN_382_0,
  output        _GEN_258_1,
  output        _GEN_304_1,
  output        _GEN_403_0,
  output        _GEN_372_0,
  output        _GEN_366_0,
  output        _GEN_267_1,
  output        _GEN_289_1,
  output        _GEN_388_0,
  output        _GEN_397_0,
  output        _GEN_252_1,
  output        _GEN_450_0,
  output        _GEN_351_0,
  output        _GEN_453_0,
  output        _GEN_447_0,
  output        _GEN_438_0,
  output        _GEN_333_0,
  output        _GEN_240_1,
  output        _GEN_339_0,
  output        _GEN_375_0,
  output        _GEN_261_1,
  output        _GEN_255_1,
  output        _GEN_360_0,
  output        _GEN_432_0,
  output        _GEN_286_1,
  output        _GEN_276_1,
  output        _GEN_459_0,
  output        _GEN_385_0,
  output        _GEN_354_0,
  output        _GEN_234_1,
  output        _GEN_3_3,
  output        _GEN_146_0,
  output        _GEN_441_0,
  output        _GEN_321_1,
  output        _GEN_348_0,
  output        _GEN_357_0,
  output        _GEN_243_1,
  output        _GEN_462_0,
  output        _GEN_456_0,
  output        _GEN_342_0,
  output        _GEN_420_0,
  output        _GEN_414_0,
  output        _GEN_336_0,
  output        _GEN_435_0,
  output        _GEN_249_1,
  output        _GEN_237_1,
  output        _GEN_315_1,
  output        _GEN_264_1,
  output        _GEN_363_0,
  output        _GEN_246_1,
  output        _GEN_150_1,
  output        _GEN_330_0,
  output        _GEN_7_3,
  output        _GEN_297_1,
  output        _GEN_345_0,
  output        _GEN_396_0,
  output        _GEN_408_0,
  output        _GEN_423_0,
  output        _GEN_309_1,
  output        _GEN_303_1,
  output        _GEN_417_0,
  output        _GEN_429_0,
  output        _GEN_444_0,
  output        _GEN_324_0,
  output        _GEN_402_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
`endif // RANDOMIZE_REG_INIT
  reg  reg_mstatus_mpie; // @[csr.scala 163:24]
  reg  reg_mstatus_mie; // @[csr.scala 163:24]
  reg [31:0] reg_mepc; // @[csr.scala 164:21]
  reg [31:0] reg_mcause; // @[csr.scala 165:23]
  reg [31:0] reg_mtval; // @[csr.scala 166:22]
  reg [31:0] reg_mscratch; // @[csr.scala 167:25]
  reg [31:0] reg_medeleg; // @[csr.scala 169:24]
  reg  reg_mip_mtip; // @[csr.scala 171:20]
  reg  reg_mip_msip; // @[csr.scala 171:20]
  reg  reg_mie_mtip; // @[csr.scala 172:20]
  reg  reg_mie_msip; // @[csr.scala 172:20]
  reg [5:0] _T_176; // @[util.scala 114:37]
  wire [6:0] _T_177 = _T_176 + 6'h1; // @[util.scala 115:33]
  reg [57:0] _T_180; // @[util.scala 119:27]
  wire [57:0] _T_184 = _T_180 + 58'h1; // @[util.scala 120:43]
  wire [63:0] _T_185 = {_T_180,_T_176}; // @[Cat.scala 30:58]
  reg [5:0] _T_188; // @[util.scala 114:37]
  wire [5:0] _GEN_153 = {{5'd0}, io_retire}; // @[util.scala 115:33]
  wire [6:0] _T_189 = _T_188 + _GEN_153; // @[util.scala 115:33]
  reg [57:0] _T_192; // @[util.scala 119:27]
  wire [57:0] _T_196 = _T_192 + 58'h1; // @[util.scala 120:43]
  wire [63:0] _T_197 = {_T_192,_T_188}; // @[Cat.scala 30:58]
  reg [39:0] _T_200; // @[util.scala 114:75]
  wire [40:0] _T_201 = {{1'd0}, _T_200}; // @[util.scala 115:33]
  reg [39:0] _T_203; // @[util.scala 114:75]
  wire [40:0] _T_204 = {{1'd0}, _T_203}; // @[util.scala 115:33]
  reg [39:0] _T_206; // @[util.scala 114:75]
  wire [40:0] _T_207 = {{1'd0}, _T_206}; // @[util.scala 115:33]
  reg [39:0] _T_209; // @[util.scala 114:75]
  wire [40:0] _T_210 = {{1'd0}, _T_209}; // @[util.scala 115:33]
  reg [39:0] _T_212; // @[util.scala 114:75]
  wire [40:0] _T_213 = {{1'd0}, _T_212}; // @[util.scala 115:33]
  reg [39:0] _T_215; // @[util.scala 114:75]
  wire [40:0] _T_216 = {{1'd0}, _T_215}; // @[util.scala 115:33]
  reg [39:0] _T_218; // @[util.scala 114:75]
  wire [40:0] _T_219 = {{1'd0}, _T_218}; // @[util.scala 115:33]
  reg [39:0] _T_221; // @[util.scala 114:75]
  wire [40:0] _T_222 = {{1'd0}, _T_221}; // @[util.scala 115:33]
  reg [39:0] _T_224; // @[util.scala 114:75]
  wire [40:0] _T_225 = {{1'd0}, _T_224}; // @[util.scala 115:33]
  reg [39:0] _T_227; // @[util.scala 114:75]
  wire [40:0] _T_228 = {{1'd0}, _T_227}; // @[util.scala 115:33]
  reg [39:0] _T_230; // @[util.scala 114:75]
  wire [40:0] _T_231 = {{1'd0}, _T_230}; // @[util.scala 115:33]
  reg [39:0] _T_233; // @[util.scala 114:75]
  wire [40:0] _T_234 = {{1'd0}, _T_233}; // @[util.scala 115:33]
  reg [39:0] _T_236; // @[util.scala 114:75]
  wire [40:0] _T_237 = {{1'd0}, _T_236}; // @[util.scala 115:33]
  reg [39:0] _T_239; // @[util.scala 114:75]
  wire [40:0] _T_240 = {{1'd0}, _T_239}; // @[util.scala 115:33]
  reg [39:0] _T_242; // @[util.scala 114:75]
  wire [40:0] _T_243 = {{1'd0}, _T_242}; // @[util.scala 115:33]
  reg [39:0] _T_245; // @[util.scala 114:75]
  wire [40:0] _T_246 = {{1'd0}, _T_245}; // @[util.scala 115:33]
  reg [39:0] _T_248; // @[util.scala 114:75]
  wire [40:0] _T_249 = {{1'd0}, _T_248}; // @[util.scala 115:33]
  reg [39:0] _T_251; // @[util.scala 114:75]
  wire [40:0] _T_252 = {{1'd0}, _T_251}; // @[util.scala 115:33]
  reg [39:0] _T_254; // @[util.scala 114:75]
  wire [40:0] _T_255 = {{1'd0}, _T_254}; // @[util.scala 115:33]
  reg [39:0] _T_257; // @[util.scala 114:75]
  wire [40:0] _T_258 = {{1'd0}, _T_257}; // @[util.scala 115:33]
  reg [39:0] _T_260; // @[util.scala 114:75]
  wire [40:0] _T_261 = {{1'd0}, _T_260}; // @[util.scala 115:33]
  reg [39:0] _T_263; // @[util.scala 114:75]
  wire [40:0] _T_264 = {{1'd0}, _T_263}; // @[util.scala 115:33]
  reg [39:0] _T_266; // @[util.scala 114:75]
  wire [40:0] _T_267 = {{1'd0}, _T_266}; // @[util.scala 115:33]
  reg [39:0] _T_269; // @[util.scala 114:75]
  wire [40:0] _T_270 = {{1'd0}, _T_269}; // @[util.scala 115:33]
  reg [39:0] _T_272; // @[util.scala 114:75]
  wire [40:0] _T_273 = {{1'd0}, _T_272}; // @[util.scala 115:33]
  reg [39:0] _T_275; // @[util.scala 114:75]
  wire [40:0] _T_276 = {{1'd0}, _T_275}; // @[util.scala 115:33]
  reg [39:0] _T_278; // @[util.scala 114:75]
  wire [40:0] _T_279 = {{1'd0}, _T_278}; // @[util.scala 115:33]
  reg [39:0] _T_281; // @[util.scala 114:75]
  wire [40:0] _T_282 = {{1'd0}, _T_281}; // @[util.scala 115:33]
  reg [39:0] _T_284; // @[util.scala 114:75]
  wire [40:0] _T_285 = {{1'd0}, _T_284}; // @[util.scala 115:33]
  reg [39:0] _T_287; // @[util.scala 114:75]
  wire [40:0] _T_288 = {{1'd0}, _T_287}; // @[util.scala 115:33]
  reg [39:0] _T_290; // @[util.scala 114:75]
  wire [40:0] _T_291 = {{1'd0}, _T_290}; // @[util.scala 115:33]
  reg [39:0] _T_293; // @[util.scala 114:75]
  wire [40:0] _T_294 = {{1'd0}, _T_293}; // @[util.scala 115:33]
  reg [31:0] reg_dpc; // @[csr.scala 188:20]
  reg [31:0] reg_dscratch; // @[csr.scala 189:25]
  reg  reg_dcsr_ebreakm; // @[csr.scala 194:21]
  reg  reg_dcsr_step; // @[csr.scala 194:21]
  wire  system_insn = io_rw_cmd == 3'h4; // @[csr.scala 196:31]
  wire  _T_410 = io_rw_cmd != 3'h0; // @[csr.scala 197:27]
  wire  _T_412 = ~system_insn; // @[csr.scala 197:39]
  wire  cpu_ren = _T_410 & _T_412; // @[csr.scala 197:36]
  wire [4:0] _T_416 = {io_status_upie,io_status_mie,io_status_hie,io_status_sie,io_status_uie};
  wire [12:0] _T_422 = {io_status_mpp,io_status_hpp,io_status_spp,io_status_mpie,io_status_hpie,io_status_spie,_T_416};
  wire [7:0] _T_427 = {io_status_tvm,io_status_mxr,io_status_sum,io_status_mprv,io_status_xs,io_status_fs};
  wire [34:0] read_mstatus = {io_status_debug,io_status_prv,io_status_sd,io_status_zero1,io_status_tsr,io_status_tw,_T_427,_T_422};
  wire [15:0] _T_454 = {8'h0,reg_mip_mtip,1'h0,2'h0,reg_mip_msip,1'h0,2'h0};
  wire [15:0] _T_469 = {8'h0,reg_mie_mtip,1'h0,2'h0,reg_mie_msip,1'h0,2'h0};
  wire [31:0] _T_483 = {4'h4,12'h0,reg_dcsr_ebreakm,4'h0,6'h0,2'h0,reg_dcsr_step,2'h3}; // @[csr.scala 222:27]
  wire  _T_487 = io_decode_csr == 12'hb00; // @[csr.scala 259:76]
  wire  _T_489 = io_decode_csr == 12'hb02; // @[csr.scala 259:76]
  wire  _T_491 = io_decode_csr == 12'hf13; // @[csr.scala 259:76]
  wire  _T_497 = io_decode_csr == 12'h301; // @[csr.scala 259:76]
  wire  _T_499 = io_decode_csr == 12'h300; // @[csr.scala 259:76]
  wire  _T_501 = io_decode_csr == 12'h305; // @[csr.scala 259:76]
  wire  _T_503 = io_decode_csr == 12'h344; // @[csr.scala 259:76]
  wire  _T_505 = io_decode_csr == 12'h304; // @[csr.scala 259:76]
  wire  _T_507 = io_decode_csr == 12'h340; // @[csr.scala 259:76]
  wire  _T_509 = io_decode_csr == 12'h341; // @[csr.scala 259:76]
  wire  _T_511 = io_decode_csr == 12'h343; // @[csr.scala 259:76]
  wire  _T_513 = io_decode_csr == 12'h342; // @[csr.scala 259:76]
  wire  _T_517 = io_decode_csr == 12'h7b0; // @[csr.scala 259:76]
  wire  _T_519 = io_decode_csr == 12'h7b1; // @[csr.scala 259:76]
  wire  _T_521 = io_decode_csr == 12'h7b2; // @[csr.scala 259:76]
  wire  _T_523 = io_decode_csr == 12'h302; // @[csr.scala 259:76]
  wire  _T_525 = io_decode_csr == 12'hb03; // @[csr.scala 259:76]
  wire  _T_527 = io_decode_csr == 12'hb83; // @[csr.scala 259:76]
  wire  _T_529 = io_decode_csr == 12'hb04; // @[csr.scala 259:76]
  wire  _T_531 = io_decode_csr == 12'hb84; // @[csr.scala 259:76]
  wire  _T_533 = io_decode_csr == 12'hb05; // @[csr.scala 259:76]
  wire  _T_535 = io_decode_csr == 12'hb85; // @[csr.scala 259:76]
  wire  _T_537 = io_decode_csr == 12'hb06; // @[csr.scala 259:76]
  wire  _T_539 = io_decode_csr == 12'hb86; // @[csr.scala 259:76]
  wire  _T_541 = io_decode_csr == 12'hb07; // @[csr.scala 259:76]
  wire  _T_543 = io_decode_csr == 12'hb87; // @[csr.scala 259:76]
  wire  _T_545 = io_decode_csr == 12'hb08; // @[csr.scala 259:76]
  wire  _T_547 = io_decode_csr == 12'hb88; // @[csr.scala 259:76]
  wire  _T_549 = io_decode_csr == 12'hb09; // @[csr.scala 259:76]
  wire  _T_551 = io_decode_csr == 12'hb89; // @[csr.scala 259:76]
  wire  _T_553 = io_decode_csr == 12'hb0a; // @[csr.scala 259:76]
  wire  _T_555 = io_decode_csr == 12'hb8a; // @[csr.scala 259:76]
  wire  _T_557 = io_decode_csr == 12'hb0b; // @[csr.scala 259:76]
  wire  _T_559 = io_decode_csr == 12'hb8b; // @[csr.scala 259:76]
  wire  _T_561 = io_decode_csr == 12'hb0c; // @[csr.scala 259:76]
  wire  _T_563 = io_decode_csr == 12'hb8c; // @[csr.scala 259:76]
  wire  _T_565 = io_decode_csr == 12'hb0d; // @[csr.scala 259:76]
  wire  _T_567 = io_decode_csr == 12'hb8d; // @[csr.scala 259:76]
  wire  _T_569 = io_decode_csr == 12'hb0e; // @[csr.scala 259:76]
  wire  _T_571 = io_decode_csr == 12'hb8e; // @[csr.scala 259:76]
  wire  _T_573 = io_decode_csr == 12'hb0f; // @[csr.scala 259:76]
  wire  _T_575 = io_decode_csr == 12'hb8f; // @[csr.scala 259:76]
  wire  _T_577 = io_decode_csr == 12'hb10; // @[csr.scala 259:76]
  wire  _T_579 = io_decode_csr == 12'hb90; // @[csr.scala 259:76]
  wire  _T_581 = io_decode_csr == 12'hb11; // @[csr.scala 259:76]
  wire  _T_583 = io_decode_csr == 12'hb91; // @[csr.scala 259:76]
  wire  _T_585 = io_decode_csr == 12'hb12; // @[csr.scala 259:76]
  wire  _T_587 = io_decode_csr == 12'hb92; // @[csr.scala 259:76]
  wire  _T_589 = io_decode_csr == 12'hb13; // @[csr.scala 259:76]
  wire  _T_591 = io_decode_csr == 12'hb93; // @[csr.scala 259:76]
  wire  _T_593 = io_decode_csr == 12'hb14; // @[csr.scala 259:76]
  wire  _T_595 = io_decode_csr == 12'hb94; // @[csr.scala 259:76]
  wire  _T_597 = io_decode_csr == 12'hb15; // @[csr.scala 259:76]
  wire  _T_599 = io_decode_csr == 12'hb95; // @[csr.scala 259:76]
  wire  _T_601 = io_decode_csr == 12'hb16; // @[csr.scala 259:76]
  wire  _T_603 = io_decode_csr == 12'hb96; // @[csr.scala 259:76]
  wire  _T_605 = io_decode_csr == 12'hb17; // @[csr.scala 259:76]
  wire  _T_607 = io_decode_csr == 12'hb97; // @[csr.scala 259:76]
  wire  _T_609 = io_decode_csr == 12'hb18; // @[csr.scala 259:76]
  wire  _T_611 = io_decode_csr == 12'hb98; // @[csr.scala 259:76]
  wire  _T_613 = io_decode_csr == 12'hb19; // @[csr.scala 259:76]
  wire  _T_615 = io_decode_csr == 12'hb99; // @[csr.scala 259:76]
  wire  _T_617 = io_decode_csr == 12'hb1a; // @[csr.scala 259:76]
  wire  _T_619 = io_decode_csr == 12'hb9a; // @[csr.scala 259:76]
  wire  _T_621 = io_decode_csr == 12'hb1b; // @[csr.scala 259:76]
  wire  _T_623 = io_decode_csr == 12'hb9b; // @[csr.scala 259:76]
  wire  _T_625 = io_decode_csr == 12'hb1c; // @[csr.scala 259:76]
  wire  _T_627 = io_decode_csr == 12'hb9c; // @[csr.scala 259:76]
  wire  _T_629 = io_decode_csr == 12'hb1d; // @[csr.scala 259:76]
  wire  _T_631 = io_decode_csr == 12'hb9d; // @[csr.scala 259:76]
  wire  _T_633 = io_decode_csr == 12'hb1e; // @[csr.scala 259:76]
  wire  _T_635 = io_decode_csr == 12'hb9e; // @[csr.scala 259:76]
  wire  _T_637 = io_decode_csr == 12'hb1f; // @[csr.scala 259:76]
  wire  _T_639 = io_decode_csr == 12'hb9f; // @[csr.scala 259:76]
  wire  _T_641 = io_decode_csr == 12'hb20; // @[csr.scala 259:76]
  wire  _T_643 = io_decode_csr == 12'hba0; // @[csr.scala 259:76]
  wire  _T_645 = io_decode_csr == 12'hb21; // @[csr.scala 259:76]
  wire  _T_647 = io_decode_csr == 12'hba1; // @[csr.scala 259:76]
  wire  _T_649 = io_decode_csr == 12'hb22; // @[csr.scala 259:76]
  wire  _T_651 = io_decode_csr == 12'hba2; // @[csr.scala 259:76]
  wire  _T_653 = io_decode_csr == 12'hb80; // @[csr.scala 259:76]
  wire  _T_655 = io_decode_csr == 12'hb82; // @[csr.scala 259:76]
  wire [1:0] _T_658 = ~io_decode_csr[11:10]; // @[csr.scala 262:40]
  wire  read_only = _T_658 == 2'h0; // @[csr.scala 262:40]
  wire  _T_660 = io_rw_cmd != 3'h5; // @[csr.scala 263:38]
  wire  cpu_wen = cpu_ren & _T_660; // @[csr.scala 263:25]
  wire  _T_663 = ~read_only; // @[csr.scala 264:24]
  wire  wen = cpu_wen & _T_663; // @[csr.scala 264:21]
  wire  _T_664 = io_rw_cmd == 3'h2; // @[util.scala 25:47]
  wire  _T_665 = io_rw_cmd == 3'h3; // @[util.scala 25:47]
  wire  _T_666 = _T_664 | _T_665; // @[util.scala 25:62]
  wire [31:0] _T_668 = _T_666 ? io_rw_rdata : 32'h0; // @[csr.scala 390:9]
  wire [31:0] _T_669 = _T_668 | io_rw_wdata; // @[csr.scala 390:53]
  wire [31:0] _T_672 = _T_665 ? io_rw_wdata : 32'h0; // @[csr.scala 390:68]
  wire [31:0] _T_673 = ~_T_672; // @[csr.scala 390:64]
  wire [31:0] wdata = _T_669 & _T_673; // @[csr.scala 390:62]
  wire [7:0] opcode = 8'h1 << io_decode_csr[2:0]; // @[csr.scala 267:20]
  wire  insn_call = system_insn & opcode[0]; // @[csr.scala 268:31]
  wire  insn_break = system_insn & opcode[1]; // @[csr.scala 269:32]
  wire  insn_ret = system_insn & opcode[2]; // @[csr.scala 270:30]
  wire  _T_962 = insn_call | insn_break; // @[csr.scala 282:24]
  wire [31:0] _GEN_4 = io_exception ? io_pc : reg_mepc; // @[csr.scala 285:23]
  wire [1:0] _T_966 = insn_ret + io_exception; // @[Bitwise.scala 48:55]
  wire  _T_968 = _T_966 <= 2'h1; // @[csr.scala 291:52]
  wire  _T_970 = _T_968 | reset; // @[csr.scala 291:9]
  wire  _T_976 = insn_ret & io_decode_csr[10]; // @[csr.scala 298:17]
  wire [31:0] _GEN_8 = _T_976 ? reg_dpc : 32'h80000004; // @[csr.scala 298:38]
  wire  _T_980 = ~io_decode_csr[10]; // @[csr.scala 305:21]
  wire  _T_981 = insn_ret & _T_980; // @[csr.scala 305:18]
  wire  _GEN_10 = _T_981 | reg_mstatus_mpie; // @[csr.scala 305:41]
  wire [31:0] _GEN_12 = _T_981 ? reg_mepc : _GEN_8; // @[csr.scala 305:41]
  wire [31:0] _GEN_13 = insn_call ? 32'h80000004 : _GEN_12; // @[csr.scala 313:18]
  wire [63:0] _T_991 = _T_487 ? _T_185 : 64'h0; // @[Mux.scala 19:72]
  wire [63:0] _T_993 = _T_489 ? _T_197 : 64'h0; // @[Mux.scala 19:72]
  wire [15:0] _T_995 = _T_491 ? 16'h8000 : 16'h0; // @[Mux.scala 19:72]
  wire [8:0] _T_1001 = _T_497 ? 9'h100 : 9'h0; // @[Mux.scala 19:72]
  wire [34:0] _T_1003 = _T_499 ? read_mstatus : 35'h0; // @[Mux.scala 19:72]
  wire [8:0] _T_1005 = _T_501 ? 9'h100 : 9'h0; // @[Mux.scala 19:72]
  wire [15:0] _T_1007 = _T_503 ? _T_454 : 16'h0; // @[Mux.scala 19:72]
  wire [15:0] _T_1009 = _T_505 ? _T_469 : 16'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1011 = _T_507 ? reg_mscratch : 32'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1013 = _T_509 ? reg_mepc : 32'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1015 = _T_511 ? reg_mtval : 32'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1017 = _T_513 ? reg_mcause : 32'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1021 = _T_517 ? _T_483 : 32'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1023 = _T_519 ? reg_dpc : 32'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1025 = _T_521 ? reg_dscratch : 32'h0; // @[Mux.scala 19:72]
  wire [31:0] _T_1027 = _T_523 ? reg_medeleg : 32'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1029 = _T_525 ? _T_200 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1031 = _T_527 ? _T_200 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1033 = _T_529 ? _T_203 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1035 = _T_531 ? _T_203 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1037 = _T_533 ? _T_206 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1039 = _T_535 ? _T_206 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1041 = _T_537 ? _T_209 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1043 = _T_539 ? _T_209 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1045 = _T_541 ? _T_212 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1047 = _T_543 ? _T_212 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1049 = _T_545 ? _T_215 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1051 = _T_547 ? _T_215 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1053 = _T_549 ? _T_218 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1055 = _T_551 ? _T_218 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1057 = _T_553 ? _T_221 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1059 = _T_555 ? _T_221 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1061 = _T_557 ? _T_224 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1063 = _T_559 ? _T_224 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1065 = _T_561 ? _T_227 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1067 = _T_563 ? _T_227 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1069 = _T_565 ? _T_230 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1071 = _T_567 ? _T_230 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1073 = _T_569 ? _T_233 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1075 = _T_571 ? _T_233 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1077 = _T_573 ? _T_236 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1079 = _T_575 ? _T_236 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1081 = _T_577 ? _T_239 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1083 = _T_579 ? _T_239 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1085 = _T_581 ? _T_242 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1087 = _T_583 ? _T_242 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1089 = _T_585 ? _T_245 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1091 = _T_587 ? _T_245 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1093 = _T_589 ? _T_248 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1095 = _T_591 ? _T_248 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1097 = _T_593 ? _T_251 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1099 = _T_595 ? _T_251 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1101 = _T_597 ? _T_254 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1103 = _T_599 ? _T_254 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1105 = _T_601 ? _T_257 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1107 = _T_603 ? _T_257 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1109 = _T_605 ? _T_260 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1111 = _T_607 ? _T_260 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1113 = _T_609 ? _T_263 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1115 = _T_611 ? _T_263 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1117 = _T_613 ? _T_266 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1119 = _T_615 ? _T_266 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1121 = _T_617 ? _T_269 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1123 = _T_619 ? _T_269 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1125 = _T_621 ? _T_272 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1127 = _T_623 ? _T_272 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1129 = _T_625 ? _T_275 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1131 = _T_627 ? _T_275 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1133 = _T_629 ? _T_278 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1135 = _T_631 ? _T_278 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1137 = _T_633 ? _T_281 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1139 = _T_635 ? _T_281 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1141 = _T_637 ? _T_284 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1143 = _T_639 ? _T_284 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1145 = _T_641 ? _T_287 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1147 = _T_643 ? _T_287 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1149 = _T_645 ? _T_290 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1151 = _T_647 ? _T_290 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1153 = _T_649 ? _T_293 : 40'h0; // @[Mux.scala 19:72]
  wire [39:0] _T_1155 = _T_651 ? _T_293 : 40'h0; // @[Mux.scala 19:72]
  wire [63:0] _T_1160 = _T_991 | _T_993; // @[Mux.scala 19:72]
  wire [63:0] _GEN_154 = {{48'd0}, _T_995}; // @[Mux.scala 19:72]
  wire [63:0] _T_1161 = _T_1160 | _GEN_154; // @[Mux.scala 19:72]
  wire [63:0] _GEN_155 = {{55'd0}, _T_1001}; // @[Mux.scala 19:72]
  wire [63:0] _T_1164 = _T_1161 | _GEN_155; // @[Mux.scala 19:72]
  wire [63:0] _GEN_156 = {{29'd0}, _T_1003}; // @[Mux.scala 19:72]
  wire [63:0] _T_1165 = _T_1164 | _GEN_156; // @[Mux.scala 19:72]
  wire [63:0] _GEN_157 = {{55'd0}, _T_1005}; // @[Mux.scala 19:72]
  wire [63:0] _T_1166 = _T_1165 | _GEN_157; // @[Mux.scala 19:72]
  wire [63:0] _GEN_158 = {{48'd0}, _T_1007}; // @[Mux.scala 19:72]
  wire [63:0] _T_1167 = _T_1166 | _GEN_158; // @[Mux.scala 19:72]
  wire [63:0] _GEN_159 = {{48'd0}, _T_1009}; // @[Mux.scala 19:72]
  wire [63:0] _T_1168 = _T_1167 | _GEN_159; // @[Mux.scala 19:72]
  wire [63:0] _GEN_160 = {{32'd0}, _T_1011}; // @[Mux.scala 19:72]
  wire [63:0] _T_1169 = _T_1168 | _GEN_160; // @[Mux.scala 19:72]
  wire [63:0] _GEN_161 = {{32'd0}, _T_1013}; // @[Mux.scala 19:72]
  wire [63:0] _T_1170 = _T_1169 | _GEN_161; // @[Mux.scala 19:72]
  wire [63:0] _GEN_162 = {{32'd0}, _T_1015}; // @[Mux.scala 19:72]
  wire [63:0] _T_1171 = _T_1170 | _GEN_162; // @[Mux.scala 19:72]
  wire [63:0] _GEN_163 = {{32'd0}, _T_1017}; // @[Mux.scala 19:72]
  wire [63:0] _T_1172 = _T_1171 | _GEN_163; // @[Mux.scala 19:72]
  wire [63:0] _GEN_164 = {{32'd0}, _T_1021}; // @[Mux.scala 19:72]
  wire [63:0] _T_1174 = _T_1172 | _GEN_164; // @[Mux.scala 19:72]
  wire [63:0] _GEN_165 = {{32'd0}, _T_1023}; // @[Mux.scala 19:72]
  wire [63:0] _T_1175 = _T_1174 | _GEN_165; // @[Mux.scala 19:72]
  wire [63:0] _GEN_166 = {{32'd0}, _T_1025}; // @[Mux.scala 19:72]
  wire [63:0] _T_1176 = _T_1175 | _GEN_166; // @[Mux.scala 19:72]
  wire [63:0] _GEN_167 = {{32'd0}, _T_1027}; // @[Mux.scala 19:72]
  wire [63:0] _T_1177 = _T_1176 | _GEN_167; // @[Mux.scala 19:72]
  wire [63:0] _GEN_168 = {{24'd0}, _T_1029}; // @[Mux.scala 19:72]
  wire [63:0] _T_1178 = _T_1177 | _GEN_168; // @[Mux.scala 19:72]
  wire [63:0] _GEN_169 = {{24'd0}, _T_1031}; // @[Mux.scala 19:72]
  wire [63:0] _T_1179 = _T_1178 | _GEN_169; // @[Mux.scala 19:72]
  wire [63:0] _GEN_170 = {{24'd0}, _T_1033}; // @[Mux.scala 19:72]
  wire [63:0] _T_1180 = _T_1179 | _GEN_170; // @[Mux.scala 19:72]
  wire [63:0] _GEN_171 = {{24'd0}, _T_1035}; // @[Mux.scala 19:72]
  wire [63:0] _T_1181 = _T_1180 | _GEN_171; // @[Mux.scala 19:72]
  wire [63:0] _GEN_172 = {{24'd0}, _T_1037}; // @[Mux.scala 19:72]
  wire [63:0] _T_1182 = _T_1181 | _GEN_172; // @[Mux.scala 19:72]
  wire [63:0] _GEN_173 = {{24'd0}, _T_1039}; // @[Mux.scala 19:72]
  wire [63:0] _T_1183 = _T_1182 | _GEN_173; // @[Mux.scala 19:72]
  wire [63:0] _GEN_174 = {{24'd0}, _T_1041}; // @[Mux.scala 19:72]
  wire [63:0] _T_1184 = _T_1183 | _GEN_174; // @[Mux.scala 19:72]
  wire [63:0] _GEN_175 = {{24'd0}, _T_1043}; // @[Mux.scala 19:72]
  wire [63:0] _T_1185 = _T_1184 | _GEN_175; // @[Mux.scala 19:72]
  wire [63:0] _GEN_176 = {{24'd0}, _T_1045}; // @[Mux.scala 19:72]
  wire [63:0] _T_1186 = _T_1185 | _GEN_176; // @[Mux.scala 19:72]
  wire [63:0] _GEN_177 = {{24'd0}, _T_1047}; // @[Mux.scala 19:72]
  wire [63:0] _T_1187 = _T_1186 | _GEN_177; // @[Mux.scala 19:72]
  wire [63:0] _GEN_178 = {{24'd0}, _T_1049}; // @[Mux.scala 19:72]
  wire [63:0] _T_1188 = _T_1187 | _GEN_178; // @[Mux.scala 19:72]
  wire [63:0] _GEN_179 = {{24'd0}, _T_1051}; // @[Mux.scala 19:72]
  wire [63:0] _T_1189 = _T_1188 | _GEN_179; // @[Mux.scala 19:72]
  wire [63:0] _GEN_180 = {{24'd0}, _T_1053}; // @[Mux.scala 19:72]
  wire [63:0] _T_1190 = _T_1189 | _GEN_180; // @[Mux.scala 19:72]
  wire [63:0] _GEN_181 = {{24'd0}, _T_1055}; // @[Mux.scala 19:72]
  wire [63:0] _T_1191 = _T_1190 | _GEN_181; // @[Mux.scala 19:72]
  wire [63:0] _GEN_182 = {{24'd0}, _T_1057}; // @[Mux.scala 19:72]
  wire [63:0] _T_1192 = _T_1191 | _GEN_182; // @[Mux.scala 19:72]
  wire [63:0] _GEN_183 = {{24'd0}, _T_1059}; // @[Mux.scala 19:72]
  wire [63:0] _T_1193 = _T_1192 | _GEN_183; // @[Mux.scala 19:72]
  wire [63:0] _GEN_184 = {{24'd0}, _T_1061}; // @[Mux.scala 19:72]
  wire [63:0] _T_1194 = _T_1193 | _GEN_184; // @[Mux.scala 19:72]
  wire [63:0] _GEN_185 = {{24'd0}, _T_1063}; // @[Mux.scala 19:72]
  wire [63:0] _T_1195 = _T_1194 | _GEN_185; // @[Mux.scala 19:72]
  wire [63:0] _GEN_186 = {{24'd0}, _T_1065}; // @[Mux.scala 19:72]
  wire [63:0] _T_1196 = _T_1195 | _GEN_186; // @[Mux.scala 19:72]
  wire [63:0] _GEN_187 = {{24'd0}, _T_1067}; // @[Mux.scala 19:72]
  wire [63:0] _T_1197 = _T_1196 | _GEN_187; // @[Mux.scala 19:72]
  wire [63:0] _GEN_188 = {{24'd0}, _T_1069}; // @[Mux.scala 19:72]
  wire [63:0] _T_1198 = _T_1197 | _GEN_188; // @[Mux.scala 19:72]
  wire [63:0] _GEN_189 = {{24'd0}, _T_1071}; // @[Mux.scala 19:72]
  wire [63:0] _T_1199 = _T_1198 | _GEN_189; // @[Mux.scala 19:72]
  wire [63:0] _GEN_190 = {{24'd0}, _T_1073}; // @[Mux.scala 19:72]
  wire [63:0] _T_1200 = _T_1199 | _GEN_190; // @[Mux.scala 19:72]
  wire [63:0] _GEN_191 = {{24'd0}, _T_1075}; // @[Mux.scala 19:72]
  wire [63:0] _T_1201 = _T_1200 | _GEN_191; // @[Mux.scala 19:72]
  wire [63:0] _GEN_192 = {{24'd0}, _T_1077}; // @[Mux.scala 19:72]
  wire [63:0] _T_1202 = _T_1201 | _GEN_192; // @[Mux.scala 19:72]
  wire [63:0] _GEN_193 = {{24'd0}, _T_1079}; // @[Mux.scala 19:72]
  wire [63:0] _T_1203 = _T_1202 | _GEN_193; // @[Mux.scala 19:72]
  wire [63:0] _GEN_194 = {{24'd0}, _T_1081}; // @[Mux.scala 19:72]
  wire [63:0] _T_1204 = _T_1203 | _GEN_194; // @[Mux.scala 19:72]
  wire [63:0] _GEN_195 = {{24'd0}, _T_1083}; // @[Mux.scala 19:72]
  wire [63:0] _T_1205 = _T_1204 | _GEN_195; // @[Mux.scala 19:72]
  wire [63:0] _GEN_196 = {{24'd0}, _T_1085}; // @[Mux.scala 19:72]
  wire [63:0] _T_1206 = _T_1205 | _GEN_196; // @[Mux.scala 19:72]
  wire [63:0] _GEN_197 = {{24'd0}, _T_1087}; // @[Mux.scala 19:72]
  wire [63:0] _T_1207 = _T_1206 | _GEN_197; // @[Mux.scala 19:72]
  wire [63:0] _GEN_198 = {{24'd0}, _T_1089}; // @[Mux.scala 19:72]
  wire [63:0] _T_1208 = _T_1207 | _GEN_198; // @[Mux.scala 19:72]
  wire [63:0] _GEN_199 = {{24'd0}, _T_1091}; // @[Mux.scala 19:72]
  wire [63:0] _T_1209 = _T_1208 | _GEN_199; // @[Mux.scala 19:72]
  wire [63:0] _GEN_200 = {{24'd0}, _T_1093}; // @[Mux.scala 19:72]
  wire [63:0] _T_1210 = _T_1209 | _GEN_200; // @[Mux.scala 19:72]
  wire [63:0] _GEN_201 = {{24'd0}, _T_1095}; // @[Mux.scala 19:72]
  wire [63:0] _T_1211 = _T_1210 | _GEN_201; // @[Mux.scala 19:72]
  wire [63:0] _GEN_202 = {{24'd0}, _T_1097}; // @[Mux.scala 19:72]
  wire [63:0] _T_1212 = _T_1211 | _GEN_202; // @[Mux.scala 19:72]
  wire [63:0] _GEN_203 = {{24'd0}, _T_1099}; // @[Mux.scala 19:72]
  wire [63:0] _T_1213 = _T_1212 | _GEN_203; // @[Mux.scala 19:72]
  wire [63:0] _GEN_204 = {{24'd0}, _T_1101}; // @[Mux.scala 19:72]
  wire [63:0] _T_1214 = _T_1213 | _GEN_204; // @[Mux.scala 19:72]
  wire [63:0] _GEN_205 = {{24'd0}, _T_1103}; // @[Mux.scala 19:72]
  wire [63:0] _T_1215 = _T_1214 | _GEN_205; // @[Mux.scala 19:72]
  wire [63:0] _GEN_206 = {{24'd0}, _T_1105}; // @[Mux.scala 19:72]
  wire [63:0] _T_1216 = _T_1215 | _GEN_206; // @[Mux.scala 19:72]
  wire [63:0] _GEN_207 = {{24'd0}, _T_1107}; // @[Mux.scala 19:72]
  wire [63:0] _T_1217 = _T_1216 | _GEN_207; // @[Mux.scala 19:72]
  wire [63:0] _GEN_208 = {{24'd0}, _T_1109}; // @[Mux.scala 19:72]
  wire [63:0] _T_1218 = _T_1217 | _GEN_208; // @[Mux.scala 19:72]
  wire [63:0] _GEN_209 = {{24'd0}, _T_1111}; // @[Mux.scala 19:72]
  wire [63:0] _T_1219 = _T_1218 | _GEN_209; // @[Mux.scala 19:72]
  wire [63:0] _GEN_210 = {{24'd0}, _T_1113}; // @[Mux.scala 19:72]
  wire [63:0] _T_1220 = _T_1219 | _GEN_210; // @[Mux.scala 19:72]
  wire [63:0] _GEN_211 = {{24'd0}, _T_1115}; // @[Mux.scala 19:72]
  wire [63:0] _T_1221 = _T_1220 | _GEN_211; // @[Mux.scala 19:72]
  wire [63:0] _GEN_212 = {{24'd0}, _T_1117}; // @[Mux.scala 19:72]
  wire [63:0] _T_1222 = _T_1221 | _GEN_212; // @[Mux.scala 19:72]
  wire [63:0] _GEN_213 = {{24'd0}, _T_1119}; // @[Mux.scala 19:72]
  wire [63:0] _T_1223 = _T_1222 | _GEN_213; // @[Mux.scala 19:72]
  wire [63:0] _GEN_214 = {{24'd0}, _T_1121}; // @[Mux.scala 19:72]
  wire [63:0] _T_1224 = _T_1223 | _GEN_214; // @[Mux.scala 19:72]
  wire [63:0] _GEN_215 = {{24'd0}, _T_1123}; // @[Mux.scala 19:72]
  wire [63:0] _T_1225 = _T_1224 | _GEN_215; // @[Mux.scala 19:72]
  wire [63:0] _GEN_216 = {{24'd0}, _T_1125}; // @[Mux.scala 19:72]
  wire [63:0] _T_1226 = _T_1225 | _GEN_216; // @[Mux.scala 19:72]
  wire [63:0] _GEN_217 = {{24'd0}, _T_1127}; // @[Mux.scala 19:72]
  wire [63:0] _T_1227 = _T_1226 | _GEN_217; // @[Mux.scala 19:72]
  wire [63:0] _GEN_218 = {{24'd0}, _T_1129}; // @[Mux.scala 19:72]
  wire [63:0] _T_1228 = _T_1227 | _GEN_218; // @[Mux.scala 19:72]
  wire [63:0] _GEN_219 = {{24'd0}, _T_1131}; // @[Mux.scala 19:72]
  wire [63:0] _T_1229 = _T_1228 | _GEN_219; // @[Mux.scala 19:72]
  wire [63:0] _GEN_220 = {{24'd0}, _T_1133}; // @[Mux.scala 19:72]
  wire [63:0] _T_1230 = _T_1229 | _GEN_220; // @[Mux.scala 19:72]
  wire [63:0] _GEN_221 = {{24'd0}, _T_1135}; // @[Mux.scala 19:72]
  wire [63:0] _T_1231 = _T_1230 | _GEN_221; // @[Mux.scala 19:72]
  wire [63:0] _GEN_222 = {{24'd0}, _T_1137}; // @[Mux.scala 19:72]
  wire [63:0] _T_1232 = _T_1231 | _GEN_222; // @[Mux.scala 19:72]
  wire [63:0] _GEN_223 = {{24'd0}, _T_1139}; // @[Mux.scala 19:72]
  wire [63:0] _T_1233 = _T_1232 | _GEN_223; // @[Mux.scala 19:72]
  wire [63:0] _GEN_224 = {{24'd0}, _T_1141}; // @[Mux.scala 19:72]
  wire [63:0] _T_1234 = _T_1233 | _GEN_224; // @[Mux.scala 19:72]
  wire [63:0] _GEN_225 = {{24'd0}, _T_1143}; // @[Mux.scala 19:72]
  wire [63:0] _T_1235 = _T_1234 | _GEN_225; // @[Mux.scala 19:72]
  wire [63:0] _GEN_226 = {{24'd0}, _T_1145}; // @[Mux.scala 19:72]
  wire [63:0] _T_1236 = _T_1235 | _GEN_226; // @[Mux.scala 19:72]
  wire [63:0] _GEN_227 = {{24'd0}, _T_1147}; // @[Mux.scala 19:72]
  wire [63:0] _T_1237 = _T_1236 | _GEN_227; // @[Mux.scala 19:72]
  wire [63:0] _GEN_228 = {{24'd0}, _T_1149}; // @[Mux.scala 19:72]
  wire [63:0] _T_1238 = _T_1237 | _GEN_228; // @[Mux.scala 19:72]
  wire [63:0] _GEN_229 = {{24'd0}, _T_1151}; // @[Mux.scala 19:72]
  wire [63:0] _T_1239 = _T_1238 | _GEN_229; // @[Mux.scala 19:72]
  wire [63:0] _GEN_230 = {{24'd0}, _T_1153}; // @[Mux.scala 19:72]
  wire [63:0] _T_1240 = _T_1239 | _GEN_230; // @[Mux.scala 19:72]
  wire [63:0] _GEN_231 = {{24'd0}, _T_1155}; // @[Mux.scala 19:72]
  wire [63:0] _T_1241 = _T_1240 | _GEN_231; // @[Mux.scala 19:72]
  wire [34:0] _T_1270 = {{3'd0}, wdata};
  wire [39:0] _T_1338 = {wdata[7:0],_T_200[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_24 = _T_527 ? {{1'd0}, _T_1338} : _T_201; // @[csr.scala 386:29]
  wire [39:0] _T_1340 = {_T_200[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_25 = _T_525 ? {{1'd0}, _T_1340} : _GEN_24; // @[csr.scala 387:29]
  wire [39:0] _T_1343 = {wdata[7:0],_T_203[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_26 = _T_531 ? {{1'd0}, _T_1343} : _T_204; // @[csr.scala 386:29]
  wire [39:0] _T_1345 = {_T_203[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_27 = _T_529 ? {{1'd0}, _T_1345} : _GEN_26; // @[csr.scala 387:29]
  wire [39:0] _T_1348 = {wdata[7:0],_T_206[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_28 = _T_535 ? {{1'd0}, _T_1348} : _T_207; // @[csr.scala 386:29]
  wire [39:0] _T_1350 = {_T_206[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_29 = _T_533 ? {{1'd0}, _T_1350} : _GEN_28; // @[csr.scala 387:29]
  wire [39:0] _T_1353 = {wdata[7:0],_T_209[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_30 = _T_539 ? {{1'd0}, _T_1353} : _T_210; // @[csr.scala 386:29]
  wire [39:0] _T_1355 = {_T_209[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_31 = _T_537 ? {{1'd0}, _T_1355} : _GEN_30; // @[csr.scala 387:29]
  wire [39:0] _T_1358 = {wdata[7:0],_T_212[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_32 = _T_543 ? {{1'd0}, _T_1358} : _T_213; // @[csr.scala 386:29]
  wire [39:0] _T_1360 = {_T_212[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_33 = _T_541 ? {{1'd0}, _T_1360} : _GEN_32; // @[csr.scala 387:29]
  wire [39:0] _T_1363 = {wdata[7:0],_T_215[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_34 = _T_547 ? {{1'd0}, _T_1363} : _T_216; // @[csr.scala 386:29]
  wire [39:0] _T_1365 = {_T_215[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_35 = _T_545 ? {{1'd0}, _T_1365} : _GEN_34; // @[csr.scala 387:29]
  wire [39:0] _T_1368 = {wdata[7:0],_T_218[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_36 = _T_551 ? {{1'd0}, _T_1368} : _T_219; // @[csr.scala 386:29]
  wire [39:0] _T_1370 = {_T_218[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_37 = _T_549 ? {{1'd0}, _T_1370} : _GEN_36; // @[csr.scala 387:29]
  wire [39:0] _T_1373 = {wdata[7:0],_T_221[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_38 = _T_555 ? {{1'd0}, _T_1373} : _T_222; // @[csr.scala 386:29]
  wire [39:0] _T_1375 = {_T_221[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_39 = _T_553 ? {{1'd0}, _T_1375} : _GEN_38; // @[csr.scala 387:29]
  wire [39:0] _T_1378 = {wdata[7:0],_T_224[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_40 = _T_559 ? {{1'd0}, _T_1378} : _T_225; // @[csr.scala 386:29]
  wire [39:0] _T_1380 = {_T_224[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_41 = _T_557 ? {{1'd0}, _T_1380} : _GEN_40; // @[csr.scala 387:29]
  wire [39:0] _T_1383 = {wdata[7:0],_T_227[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_42 = _T_563 ? {{1'd0}, _T_1383} : _T_228; // @[csr.scala 386:29]
  wire [39:0] _T_1385 = {_T_227[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_43 = _T_561 ? {{1'd0}, _T_1385} : _GEN_42; // @[csr.scala 387:29]
  wire [39:0] _T_1388 = {wdata[7:0],_T_230[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_44 = _T_567 ? {{1'd0}, _T_1388} : _T_231; // @[csr.scala 386:29]
  wire [39:0] _T_1390 = {_T_230[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_45 = _T_565 ? {{1'd0}, _T_1390} : _GEN_44; // @[csr.scala 387:29]
  wire [39:0] _T_1393 = {wdata[7:0],_T_233[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_46 = _T_571 ? {{1'd0}, _T_1393} : _T_234; // @[csr.scala 386:29]
  wire [39:0] _T_1395 = {_T_233[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_47 = _T_569 ? {{1'd0}, _T_1395} : _GEN_46; // @[csr.scala 387:29]
  wire [39:0] _T_1398 = {wdata[7:0],_T_236[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_48 = _T_575 ? {{1'd0}, _T_1398} : _T_237; // @[csr.scala 386:29]
  wire [39:0] _T_1400 = {_T_236[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_49 = _T_573 ? {{1'd0}, _T_1400} : _GEN_48; // @[csr.scala 387:29]
  wire [39:0] _T_1403 = {wdata[7:0],_T_239[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_50 = _T_579 ? {{1'd0}, _T_1403} : _T_240; // @[csr.scala 386:29]
  wire [39:0] _T_1405 = {_T_239[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_51 = _T_577 ? {{1'd0}, _T_1405} : _GEN_50; // @[csr.scala 387:29]
  wire [39:0] _T_1408 = {wdata[7:0],_T_242[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_52 = _T_583 ? {{1'd0}, _T_1408} : _T_243; // @[csr.scala 386:29]
  wire [39:0] _T_1410 = {_T_242[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_53 = _T_581 ? {{1'd0}, _T_1410} : _GEN_52; // @[csr.scala 387:29]
  wire [39:0] _T_1413 = {wdata[7:0],_T_245[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_54 = _T_587 ? {{1'd0}, _T_1413} : _T_246; // @[csr.scala 386:29]
  wire [39:0] _T_1415 = {_T_245[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_55 = _T_585 ? {{1'd0}, _T_1415} : _GEN_54; // @[csr.scala 387:29]
  wire [39:0] _T_1418 = {wdata[7:0],_T_248[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_56 = _T_591 ? {{1'd0}, _T_1418} : _T_249; // @[csr.scala 386:29]
  wire [39:0] _T_1420 = {_T_248[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_57 = _T_589 ? {{1'd0}, _T_1420} : _GEN_56; // @[csr.scala 387:29]
  wire [39:0] _T_1423 = {wdata[7:0],_T_251[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_58 = _T_595 ? {{1'd0}, _T_1423} : _T_252; // @[csr.scala 386:29]
  wire [39:0] _T_1425 = {_T_251[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_59 = _T_593 ? {{1'd0}, _T_1425} : _GEN_58; // @[csr.scala 387:29]
  wire [39:0] _T_1428 = {wdata[7:0],_T_254[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_60 = _T_599 ? {{1'd0}, _T_1428} : _T_255; // @[csr.scala 386:29]
  wire [39:0] _T_1430 = {_T_254[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_61 = _T_597 ? {{1'd0}, _T_1430} : _GEN_60; // @[csr.scala 387:29]
  wire [39:0] _T_1433 = {wdata[7:0],_T_257[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_62 = _T_603 ? {{1'd0}, _T_1433} : _T_258; // @[csr.scala 386:29]
  wire [39:0] _T_1435 = {_T_257[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_63 = _T_601 ? {{1'd0}, _T_1435} : _GEN_62; // @[csr.scala 387:29]
  wire [39:0] _T_1438 = {wdata[7:0],_T_260[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_64 = _T_607 ? {{1'd0}, _T_1438} : _T_261; // @[csr.scala 386:29]
  wire [39:0] _T_1440 = {_T_260[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_65 = _T_605 ? {{1'd0}, _T_1440} : _GEN_64; // @[csr.scala 387:29]
  wire [39:0] _T_1443 = {wdata[7:0],_T_263[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_66 = _T_611 ? {{1'd0}, _T_1443} : _T_264; // @[csr.scala 386:29]
  wire [39:0] _T_1445 = {_T_263[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_67 = _T_609 ? {{1'd0}, _T_1445} : _GEN_66; // @[csr.scala 387:29]
  wire [39:0] _T_1448 = {wdata[7:0],_T_266[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_68 = _T_615 ? {{1'd0}, _T_1448} : _T_267; // @[csr.scala 386:29]
  wire [39:0] _T_1450 = {_T_266[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_69 = _T_613 ? {{1'd0}, _T_1450} : _GEN_68; // @[csr.scala 387:29]
  wire [39:0] _T_1453 = {wdata[7:0],_T_269[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_70 = _T_619 ? {{1'd0}, _T_1453} : _T_270; // @[csr.scala 386:29]
  wire [39:0] _T_1455 = {_T_269[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_71 = _T_617 ? {{1'd0}, _T_1455} : _GEN_70; // @[csr.scala 387:29]
  wire [39:0] _T_1458 = {wdata[7:0],_T_272[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_72 = _T_623 ? {{1'd0}, _T_1458} : _T_273; // @[csr.scala 386:29]
  wire [39:0] _T_1460 = {_T_272[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_73 = _T_621 ? {{1'd0}, _T_1460} : _GEN_72; // @[csr.scala 387:29]
  wire [39:0] _T_1463 = {wdata[7:0],_T_275[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_74 = _T_627 ? {{1'd0}, _T_1463} : _T_276; // @[csr.scala 386:29]
  wire [39:0] _T_1465 = {_T_275[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_75 = _T_625 ? {{1'd0}, _T_1465} : _GEN_74; // @[csr.scala 387:29]
  wire [39:0] _T_1468 = {wdata[7:0],_T_278[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_76 = _T_631 ? {{1'd0}, _T_1468} : _T_279; // @[csr.scala 386:29]
  wire [39:0] _T_1470 = {_T_278[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_77 = _T_629 ? {{1'd0}, _T_1470} : _GEN_76; // @[csr.scala 387:29]
  wire [39:0] _T_1473 = {wdata[7:0],_T_281[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_78 = _T_635 ? {{1'd0}, _T_1473} : _T_282; // @[csr.scala 386:29]
  wire [39:0] _T_1475 = {_T_281[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_79 = _T_633 ? {{1'd0}, _T_1475} : _GEN_78; // @[csr.scala 387:29]
  wire [39:0] _T_1478 = {wdata[7:0],_T_284[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_80 = _T_639 ? {{1'd0}, _T_1478} : _T_285; // @[csr.scala 386:29]
  wire [39:0] _T_1480 = {_T_284[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_81 = _T_637 ? {{1'd0}, _T_1480} : _GEN_80; // @[csr.scala 387:29]
  wire [39:0] _T_1483 = {wdata[7:0],_T_287[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_82 = _T_643 ? {{1'd0}, _T_1483} : _T_288; // @[csr.scala 386:29]
  wire [39:0] _T_1485 = {_T_287[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_83 = _T_641 ? {{1'd0}, _T_1485} : _GEN_82; // @[csr.scala 387:29]
  wire [39:0] _T_1488 = {wdata[7:0],_T_290[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_84 = _T_647 ? {{1'd0}, _T_1488} : _T_291; // @[csr.scala 386:29]
  wire [39:0] _T_1490 = {_T_290[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_85 = _T_645 ? {{1'd0}, _T_1490} : _GEN_84; // @[csr.scala 387:29]
  wire [39:0] _T_1493 = {wdata[7:0],_T_293[31:0]}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_86 = _T_651 ? {{1'd0}, _T_1493} : _T_294; // @[csr.scala 386:29]
  wire [39:0] _T_1495 = {_T_293[39:32],wdata}; // @[Cat.scala 30:58]
  wire [40:0] _GEN_87 = _T_649 ? {{1'd0}, _T_1495} : _GEN_86; // @[csr.scala 387:29]
  wire [63:0] _T_1498 = {wdata,_T_185[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_88 = _T_653 ? _T_1498 : {{57'd0}, _T_177}; // @[csr.scala 386:29]
  wire [63:0] _T_1501 = {_T_185[63:32],wdata}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_90 = _T_487 ? _T_1501 : _GEN_88; // @[csr.scala 387:29]
  wire [63:0] _T_1505 = {wdata,_T_197[31:0]}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_92 = _T_655 ? _T_1505 : {{57'd0}, _T_189}; // @[csr.scala 386:29]
  wire [63:0] _T_1508 = {_T_197[63:32],wdata}; // @[Cat.scala 30:58]
  wire [63:0] _GEN_94 = _T_489 ? _T_1508 : _GEN_92; // @[csr.scala 387:29]
  wire [31:0] _T_1512 = {{2'd0}, wdata[31:2]}; // @[csr.scala 368:78]
  wire [33:0] _GEN_233 = {_T_1512, 2'h0}; // @[csr.scala 368:86]
  wire [34:0] _T_1514 = {{1'd0}, _GEN_233}; // @[csr.scala 368:86]
  wire [34:0] _GEN_98 = _T_509 ? _T_1514 : {{3'd0}, _GEN_4}; // @[csr.scala 368:40]
  wire [31:0] _T_1516 = wdata & 32'h8000001f; // @[csr.scala 370:62]
  wire [40:0] _GEN_110 = wen ? _GEN_25 : _T_201; // @[csr.scala 331:14]
  wire [40:0] _GEN_111 = wen ? _GEN_27 : _T_204; // @[csr.scala 331:14]
  wire [40:0] _GEN_112 = wen ? _GEN_29 : _T_207; // @[csr.scala 331:14]
  wire [40:0] _GEN_113 = wen ? _GEN_31 : _T_210; // @[csr.scala 331:14]
  wire [40:0] _GEN_114 = wen ? _GEN_33 : _T_213; // @[csr.scala 331:14]
  wire [40:0] _GEN_115 = wen ? _GEN_35 : _T_216; // @[csr.scala 331:14]
  wire [40:0] _GEN_116 = wen ? _GEN_37 : _T_219; // @[csr.scala 331:14]
  wire [40:0] _GEN_117 = wen ? _GEN_39 : _T_222; // @[csr.scala 331:14]
  wire [40:0] _GEN_118 = wen ? _GEN_41 : _T_225; // @[csr.scala 331:14]
  wire [40:0] _GEN_119 = wen ? _GEN_43 : _T_228; // @[csr.scala 331:14]
  wire [40:0] _GEN_120 = wen ? _GEN_45 : _T_231; // @[csr.scala 331:14]
  wire [40:0] _GEN_121 = wen ? _GEN_47 : _T_234; // @[csr.scala 331:14]
  wire [40:0] _GEN_122 = wen ? _GEN_49 : _T_237; // @[csr.scala 331:14]
  wire [40:0] _GEN_123 = wen ? _GEN_51 : _T_240; // @[csr.scala 331:14]
  wire [40:0] _GEN_124 = wen ? _GEN_53 : _T_243; // @[csr.scala 331:14]
  wire [40:0] _GEN_125 = wen ? _GEN_55 : _T_246; // @[csr.scala 331:14]
  wire [40:0] _GEN_126 = wen ? _GEN_57 : _T_249; // @[csr.scala 331:14]
  wire [40:0] _GEN_127 = wen ? _GEN_59 : _T_252; // @[csr.scala 331:14]
  wire [40:0] _GEN_128 = wen ? _GEN_61 : _T_255; // @[csr.scala 331:14]
  wire [40:0] _GEN_129 = wen ? _GEN_63 : _T_258; // @[csr.scala 331:14]
  wire [40:0] _GEN_130 = wen ? _GEN_65 : _T_261; // @[csr.scala 331:14]
  wire [40:0] _GEN_131 = wen ? _GEN_67 : _T_264; // @[csr.scala 331:14]
  wire [40:0] _GEN_132 = wen ? _GEN_69 : _T_267; // @[csr.scala 331:14]
  wire [40:0] _GEN_133 = wen ? _GEN_71 : _T_270; // @[csr.scala 331:14]
  wire [40:0] _GEN_134 = wen ? _GEN_73 : _T_273; // @[csr.scala 331:14]
  wire [40:0] _GEN_135 = wen ? _GEN_75 : _T_276; // @[csr.scala 331:14]
  wire [40:0] _GEN_136 = wen ? _GEN_77 : _T_279; // @[csr.scala 331:14]
  wire [40:0] _GEN_137 = wen ? _GEN_79 : _T_282; // @[csr.scala 331:14]
  wire [40:0] _GEN_138 = wen ? _GEN_81 : _T_285; // @[csr.scala 331:14]
  wire [40:0] _GEN_139 = wen ? _GEN_83 : _T_288; // @[csr.scala 331:14]
  wire [40:0] _GEN_140 = wen ? _GEN_85 : _T_291; // @[csr.scala 331:14]
  wire [40:0] _GEN_141 = wen ? _GEN_87 : _T_294; // @[csr.scala 331:14]
  wire [63:0] _GEN_142 = wen ? _GEN_90 : {{57'd0}, _T_177}; // @[csr.scala 331:14]
  wire [63:0] _GEN_144 = wen ? _GEN_94 : {{57'd0}, _T_189}; // @[csr.scala 331:14]
  wire [34:0] _GEN_148 = wen ? _GEN_98 : {{3'd0}, _GEN_4}; // @[csr.scala 331:14]
  assign io_rw_rdata = _T_1241[31:0]; // @[csr.scala 329:15]
  assign io_eret = _T_962 | insn_ret; // @[csr.scala 282:11]
  assign io_status_debug = 1'h0; // @[csr.scala 280:13]
  assign io_status_prv = 2'h3; // @[csr.scala 280:13]
  assign io_status_sd = 1'h0; // @[csr.scala 280:13]
  assign io_status_zero1 = 8'h0; // @[csr.scala 280:13]
  assign io_status_tsr = 1'h0; // @[csr.scala 280:13]
  assign io_status_tw = 1'h0; // @[csr.scala 280:13]
  assign io_status_tvm = 1'h0; // @[csr.scala 280:13]
  assign io_status_mxr = 1'h0; // @[csr.scala 280:13]
  assign io_status_sum = 1'h0; // @[csr.scala 280:13]
  assign io_status_mprv = 1'h0; // @[csr.scala 280:13]
  assign io_status_xs = 2'h0; // @[csr.scala 280:13]
  assign io_status_fs = 2'h0; // @[csr.scala 280:13]
  assign io_status_mpp = 2'h3; // @[csr.scala 280:13]
  assign io_status_hpp = 2'h0; // @[csr.scala 280:13]
  assign io_status_spp = 1'h0; // @[csr.scala 280:13]
  assign io_status_mpie = reg_mstatus_mpie; // @[csr.scala 280:13]
  assign io_status_hpie = 1'h0; // @[csr.scala 280:13]
  assign io_status_spie = 1'h0; // @[csr.scala 280:13]
  assign io_status_upie = 1'h0; // @[csr.scala 280:13]
  assign io_status_mie = reg_mstatus_mie; // @[csr.scala 280:13]
  assign io_status_hie = 1'h0; // @[csr.scala 280:13]
  assign io_status_sie = 1'h0; // @[csr.scala 280:13]
  assign io_status_uie = 1'h0; // @[csr.scala 280:13]
  assign io_evec = insn_break ? 32'h80000004 : _GEN_13; // @[csr.scala 287:13 csr.scala 301:13 csr.scala 309:13 csr.scala 314:13 csr.scala 320:13]
  assign _GEN_411_0 = cpu_wen & _T_663;
  assign _GEN_405_0 = cpu_wen & _T_663;
  assign _GEN_426_0 = cpu_wen & _T_663;
  assign _GEN_291_0 = io_decode_csr == 12'hb97;
  assign _GEN_306_0 = io_decode_csr == 12'hb1f;
  assign _GEN_384_0 = io_decode_csr == 12'hb22;
  assign _GEN_327_0 = io_decode_csr == 12'hb86;
  assign _GEN_390_0 = io_decode_csr == 12'hb82;
  assign _GEN_285_0 = io_decode_csr == 12'hb94;
  assign _GEN_318_0 = io_decode_csr == 12'h344;
  assign _GEN_312_0 = io_decode_csr == 12'hb22;
  assign _GEN_399_0 = io_decode_csr == 12'h302;
  assign _GEN_387_0 = io_decode_csr == 12'hb00;
  assign _GEN_300_0 = io_decode_csr == 12'hb1c;
  assign _GEN_279_0 = io_decode_csr == 12'hb91;
  assign _GEN_269_0 = io_decode_csr == 12'hb8c;
  assign _GEN_378_0 = io_decode_csr == 12'hb1f;
  assign _GEN_368_0 = io_decode_csr == 12'hb1a;
  assign _GEN_377_0 = io_decode_csr == 12'hb9f;
  assign _GEN_294_0 = io_decode_csr == 12'hb19;
  assign _GEN_393_0 = io_decode_csr == 12'h7b1;
  assign _GEN_362_0 = io_decode_csr == 12'hb17;
  assign _GEN_461_0 = reset;
  assign _GEN_263_0 = io_decode_csr == 12'hb89;
  assign _GEN_449_0 = cpu_wen & _T_663;
  assign _GEN_288_0 = io_decode_csr == 12'hb16;
  assign _GEN_245_0 = io_decode_csr == 12'h342;
  assign _GEN_272_0 = io_decode_csr == 12'hb0e;
  assign _GEN_381_0 = io_decode_csr == 12'hba1;
  assign _GEN_371_0 = io_decode_csr == 12'hb9c;
  assign _GEN_266_0 = io_decode_csr == 12'hb0b;
  assign _GEN_344_0 = io_decode_csr == 12'hb0e;
  assign _GEN_282_0 = io_decode_csr == 12'hb13;
  assign _GEN_443_0 = cpu_wen & _T_663;
  assign _GEN_251_0 = io_decode_csr == 12'hb83;
  assign _GEN_350_0 = io_decode_csr == 12'hb11;
  assign _GEN_365_0 = io_decode_csr == 12'hb99;
  assign _GEN_15_0 = io_exception;
  assign _GEN_152_0 = system_insn & opcode[1];
  assign _GEN_446_0 = reset;
  assign _GEN_332_0 = io_decode_csr == 12'hb08;
  assign _GEN_326_0 = io_decode_csr == 12'hb05;
  assign _GEN_359_0 = io_decode_csr == 12'hb96;
  assign _GEN_458_0 = reset;
  assign _GEN_452_0 = reset;
  assign _GEN_347_0 = io_decode_csr == 12'hb90;
  assign _GEN_425_0 = cpu_wen & _T_663;
  assign _GEN_239_0 = io_decode_csr == 12'h305;
  assign _GEN_431_0 = cpu_wen & _T_663;
  assign _GEN_254_0 = io_decode_csr == 12'hb05;
  assign _GEN_353_0 = io_decode_csr == 12'hb93;
  assign _GEN_260_0 = io_decode_csr == 12'hb08;
  assign _GEN_275_0 = io_decode_csr == 12'hb8f;
  assign _GEN_338_0 = io_decode_csr == 12'hb0b;
  assign _GEN_374_0 = io_decode_csr == 12'hb1d;
  assign _GEN_242_0 = io_decode_csr == 12'h340;
  assign _GEN_455_0 = reset;
  assign _GEN_413_0 = cpu_wen & _T_663;
  assign _GEN_236_0 = io_decode_csr == 12'hf13;
  assign _GEN_335_0 = io_decode_csr == 12'hb8a;
  assign _GEN_434_0 = cpu_wen & _T_663;
  assign _GEN_248_1 = io_decode_csr == 12'h7b2;
  assign _GEN_257_0 = io_decode_csr == 12'hb86;
  assign _GEN_320_1 = io_decode_csr == 12'h304;
  assign _GEN_356_0 = io_decode_csr == 12'hb14;
  assign _GEN_419_0 = cpu_wen & _T_663;
  assign _GEN_314_1 = io_decode_csr == 12'h7b0;
  assign _GEN_341_0 = io_decode_csr == 12'hb8d;
  assign _GEN_440_0 = cpu_wen & _T_663;
  assign _GEN_299_1 = io_decode_csr == 12'hb9b;
  assign _GEN_398_0 = io_decode_csr == 12'h343;
  assign _GEN_407_0 = cpu_wen & _T_663;
  assign _GEN_149_1 = insn_ret & _T_980;
  assign _GEN_416_0 = cpu_wen & _T_663;
  assign _GEN_281_0 = io_decode_csr == 12'hb92;
  assign _GEN_380_0 = io_decode_csr == 12'hb20;
  assign _GEN_296_1 = io_decode_csr == 12'hb1a;
  assign _GEN_422_0 = cpu_wen & _T_663;
  assign _GEN_329_0 = io_decode_csr == 12'hb87;
  assign _GEN_6_1 = _T_664 | _T_665;
  assign _GEN_437_0 = cpu_wen & _T_663;
  assign _GEN_302_1 = io_decode_csr == 12'hb1d;
  assign _GEN_401_0 = cpu_wen & _T_663;
  assign _GEN_395_0 = io_decode_csr == 12'h341;
  assign _GEN_428_0 = cpu_wen & _T_663;
  assign _GEN_308_1 = io_decode_csr == 12'hb20;
  assign _GEN_323_0 = io_decode_csr == 12'hb84;
  assign _GEN_317_0 = io_decode_csr == 12'h300;
  assign _GEN_404_0 = cpu_wen & _T_663;
  assign _GEN_290_0 = io_decode_csr == 12'hb17;
  assign _GEN_367_0 = io_decode_csr == 12'hb9a;
  assign _GEN_284_0 = io_decode_csr == 12'hb14;
  assign _GEN_274_1 = io_decode_csr == 12'hb0f;
  assign _GEN_383_0 = io_decode_csr == 12'hba2;
  assign _GEN_373_0 = io_decode_csr == 12'hb9d;
  assign _GEN_410_0 = cpu_wen & _T_663;
  assign _GEN_305_1 = io_decode_csr == 12'hb9e;
  assign _GEN_311_1 = io_decode_csr == 12'hba1;
  assign _GEN_389_0 = io_decode_csr == 12'hb82;
  assign _GEN_268_1 = io_decode_csr == 12'hb0c;
  assign _GEN_376_0 = io_decode_csr == 12'hb1e;
  assign _GEN_454_0 = reset;
  assign _GEN_293_1 = io_decode_csr == 12'hb98;
  assign _GEN_392_0 = io_decode_csr == 12'hb02;
  assign _GEN_361_0 = io_decode_csr == 12'hb97;
  assign _GEN_287_0 = io_decode_csr == 12'hb95;
  assign _GEN_256_1 = io_decode_csr == 12'hb06;
  assign _GEN_460_0 = cpu_wen & _T_663;
  assign _GEN_278_0 = io_decode_csr == 12'hb11;
  assign _GEN_355_0 = io_decode_csr == 12'hb94;
  assign _GEN_386_0 = io_decode_csr == 12'hb80;
  assign _GEN_277_1 = io_decode_csr == 12'hb90;
  assign _GEN_262_1 = io_decode_csr == 12'hb09;
  assign _GEN_244_1 = io_decode_csr == 12'h343;
  assign _GEN_448_0 = cpu_wen & _T_663;
  assign _GEN_442_0 = cpu_wen & _T_663;
  assign _GEN_457_0 = reset;
  assign _GEN_337_0 = io_decode_csr == 12'hb8b;
  assign _GEN_364_0 = io_decode_csr == 12'hb18;
  assign _GEN_328_0 = io_decode_csr == 12'hb06;
  assign _GEN_463_0 = ~_T_970;
  assign _GEN_436_0 = cpu_wen & _T_663;
  assign _GEN_370_0 = io_decode_csr == 12'hb1b;
  assign _GEN_250_1 = io_decode_csr == 12'hb03;
  assign _GEN_265_1 = io_decode_csr == 12'hb8a;
  assign _GEN_271_1 = io_decode_csr == 12'hb8d;
  assign _GEN_349_0 = io_decode_csr == 12'hb91;
  assign _GEN_343_0 = io_decode_csr == 12'hb8e;
  assign _GEN_147_0 = insn_ret & _T_980;
  assign _GEN_352_0 = io_decode_csr == 12'hb12;
  assign _GEN_247_1 = io_decode_csr == 12'h7b1;
  assign _GEN_325_0 = io_decode_csr == 12'hb85;
  assign _GEN_151_1 = system_insn & opcode[0];
  assign _GEN_238_1 = io_decode_csr == 12'h300;
  assign _GEN_451_0 = reset;
  assign _GEN_346_0 = io_decode_csr == 12'hb0f;
  assign _GEN_409_0 = cpu_wen & _T_663;
  assign _GEN_253_1 = io_decode_csr == 12'hb84;
  assign _GEN_331_0 = io_decode_csr == 12'hb88;
  assign _GEN_11_1 = io_exception;
  assign _GEN_430_0 = cpu_wen & _T_663;
  assign _GEN_424_0 = cpu_wen & _T_663;
  assign _GEN_445_0 = reset;
  assign _GEN_310_1 = io_decode_csr == 12'hb21;
  assign _GEN_259_1 = io_decode_csr == 12'hb87;
  assign _GEN_358_0 = io_decode_csr == 12'hb15;
  assign _GEN_334_0 = io_decode_csr == 12'hb09;
  assign _GEN_412_0 = cpu_wen & _T_663;
  assign _GEN_418_0 = cpu_wen & _T_663;
  assign _GEN_427_0 = cpu_wen & _T_663;
  assign _GEN_313_1 = io_decode_csr == 12'hba2;
  assign _GEN_292_1 = io_decode_csr == 12'hb18;
  assign _GEN_241_1 = io_decode_csr == 12'h304;
  assign _GEN_340_0 = io_decode_csr == 12'hb0c;
  assign _GEN_235_1 = io_decode_csr == 12'hb02;
  assign _GEN_439_0 = cpu_wen & _T_663;
  assign _GEN_298_1 = io_decode_csr == 12'hb1b;
  assign _GEN_307_1 = io_decode_csr == 12'hb9f;
  assign _GEN_406_0 = cpu_wen & _T_663;
  assign _GEN_433_0 = cpu_wen & _T_663;
  assign _GEN_319_1 = io_decode_csr == 12'h304;
  assign _GEN_391_0 = io_decode_csr == 12'hb02;
  assign _GEN_400_0 = cpu_wen & _T_663;
  assign _GEN_415_0 = cpu_wen & _T_663;
  assign _GEN_295_1 = io_decode_csr == 12'hb99;
  assign _GEN_270_1 = io_decode_csr == 12'hb0d;
  assign _GEN_322_1 = io_decode_csr == 12'hb03;
  assign _GEN_421_0 = cpu_wen & _T_663;
  assign _GEN_280_1 = io_decode_csr == 12'hb12;
  assign _GEN_379_0 = io_decode_csr == 12'hba0;
  assign _GEN_394_0 = io_decode_csr == 12'h7b2;
  assign _GEN_369_0 = io_decode_csr == 12'hb9b;
  assign _GEN_5_2 = _T_189[6];
  assign _GEN_316_1 = io_decode_csr == 12'h300;
  assign _GEN_301_1 = io_decode_csr == 12'hb9c;
  assign _GEN_283_1 = io_decode_csr == 12'hb93;
  assign _GEN_273_1 = io_decode_csr == 12'hb8e;
  assign _GEN_382_0 = io_decode_csr == 12'hb21;
  assign _GEN_258_1 = io_decode_csr == 12'hb07;
  assign _GEN_304_1 = io_decode_csr == 12'hb1e;
  assign _GEN_403_0 = cpu_wen & _T_663;
  assign _GEN_372_0 = io_decode_csr == 12'hb1c;
  assign _GEN_366_0 = io_decode_csr == 12'hb19;
  assign _GEN_267_1 = io_decode_csr == 12'hb8b;
  assign _GEN_289_1 = io_decode_csr == 12'hb96;
  assign _GEN_388_0 = io_decode_csr == 12'hb00;
  assign _GEN_397_0 = io_decode_csr == 12'h342;
  assign _GEN_252_1 = io_decode_csr == 12'hb04;
  assign _GEN_450_0 = cpu_wen & _T_663;
  assign _GEN_351_0 = io_decode_csr == 12'hb92;
  assign _GEN_453_0 = reset;
  assign _GEN_447_0 = cpu_wen & _T_663;
  assign _GEN_438_0 = cpu_wen & _T_663;
  assign _GEN_333_0 = io_decode_csr == 12'hb89;
  assign _GEN_240_1 = io_decode_csr == 12'h344;
  assign _GEN_339_0 = io_decode_csr == 12'hb8c;
  assign _GEN_375_0 = io_decode_csr == 12'hb9e;
  assign _GEN_261_1 = io_decode_csr == 12'hb88;
  assign _GEN_255_1 = io_decode_csr == 12'hb85;
  assign _GEN_360_0 = io_decode_csr == 12'hb16;
  assign _GEN_432_0 = cpu_wen & _T_663;
  assign _GEN_286_1 = io_decode_csr == 12'hb15;
  assign _GEN_276_1 = io_decode_csr == 12'hb10;
  assign _GEN_459_0 = cpu_wen & _T_663;
  assign _GEN_385_0 = io_decode_csr == 12'hb80;
  assign _GEN_354_0 = io_decode_csr == 12'hb13;
  assign _GEN_234_1 = io_decode_csr == 12'hb00;
  assign _GEN_3_3 = _T_177[6];
  assign _GEN_146_0 = insn_ret & io_decode_csr[10];
  assign _GEN_441_0 = cpu_wen & _T_663;
  assign _GEN_321_1 = io_decode_csr == 12'hb83;
  assign _GEN_348_0 = io_decode_csr == 12'hb10;
  assign _GEN_357_0 = io_decode_csr == 12'hb95;
  assign _GEN_243_1 = io_decode_csr == 12'h341;
  assign _GEN_462_0 = reset;
  assign _GEN_456_0 = reset;
  assign _GEN_342_0 = io_decode_csr == 12'hb0d;
  assign _GEN_420_0 = cpu_wen & _T_663;
  assign _GEN_414_0 = cpu_wen & _T_663;
  assign _GEN_336_0 = io_decode_csr == 12'hb0a;
  assign _GEN_435_0 = cpu_wen & _T_663;
  assign _GEN_249_1 = io_decode_csr == 12'h302;
  assign _GEN_237_1 = io_decode_csr == 12'h301;
  assign _GEN_315_1 = io_decode_csr == 12'h7b0;
  assign _GEN_264_1 = io_decode_csr == 12'hb0a;
  assign _GEN_363_0 = io_decode_csr == 12'hb98;
  assign _GEN_246_1 = io_decode_csr == 12'h7b0;
  assign _GEN_150_1 = system_insn & opcode[0];
  assign _GEN_330_0 = io_decode_csr == 12'hb07;
  assign _GEN_7_3 = io_rw_cmd == 3'h3;
  assign _GEN_297_1 = io_decode_csr == 12'hb9a;
  assign _GEN_345_0 = io_decode_csr == 12'hb8f;
  assign _GEN_396_0 = io_decode_csr == 12'h340;
  assign _GEN_408_0 = cpu_wen & _T_663;
  assign _GEN_423_0 = cpu_wen & _T_663;
  assign _GEN_309_1 = io_decode_csr == 12'hba0;
  assign _GEN_303_1 = io_decode_csr == 12'hb9d;
  assign _GEN_417_0 = cpu_wen & _T_663;
  assign _GEN_429_0 = cpu_wen & _T_663;
  assign _GEN_444_0 = system_insn & opcode[1];
  assign _GEN_324_0 = io_decode_csr == 12'hb04;
  assign _GEN_402_0 = cpu_wen & _T_663;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mstatus_mpie = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  reg_mstatus_mie = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  reg_mepc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  reg_mcause = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_mtval = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_mscratch = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_medeleg = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_mip_mtip = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  reg_mip_msip = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  reg_mie_mtip = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  reg_mie_msip = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_176 = _RAND_11[5:0];
  _RAND_12 = {2{`RANDOM}};
  _T_180 = _RAND_12[57:0];
  _RAND_13 = {1{`RANDOM}};
  _T_188 = _RAND_13[5:0];
  _RAND_14 = {2{`RANDOM}};
  _T_192 = _RAND_14[57:0];
  _RAND_15 = {2{`RANDOM}};
  _T_200 = _RAND_15[39:0];
  _RAND_16 = {2{`RANDOM}};
  _T_203 = _RAND_16[39:0];
  _RAND_17 = {2{`RANDOM}};
  _T_206 = _RAND_17[39:0];
  _RAND_18 = {2{`RANDOM}};
  _T_209 = _RAND_18[39:0];
  _RAND_19 = {2{`RANDOM}};
  _T_212 = _RAND_19[39:0];
  _RAND_20 = {2{`RANDOM}};
  _T_215 = _RAND_20[39:0];
  _RAND_21 = {2{`RANDOM}};
  _T_218 = _RAND_21[39:0];
  _RAND_22 = {2{`RANDOM}};
  _T_221 = _RAND_22[39:0];
  _RAND_23 = {2{`RANDOM}};
  _T_224 = _RAND_23[39:0];
  _RAND_24 = {2{`RANDOM}};
  _T_227 = _RAND_24[39:0];
  _RAND_25 = {2{`RANDOM}};
  _T_230 = _RAND_25[39:0];
  _RAND_26 = {2{`RANDOM}};
  _T_233 = _RAND_26[39:0];
  _RAND_27 = {2{`RANDOM}};
  _T_236 = _RAND_27[39:0];
  _RAND_28 = {2{`RANDOM}};
  _T_239 = _RAND_28[39:0];
  _RAND_29 = {2{`RANDOM}};
  _T_242 = _RAND_29[39:0];
  _RAND_30 = {2{`RANDOM}};
  _T_245 = _RAND_30[39:0];
  _RAND_31 = {2{`RANDOM}};
  _T_248 = _RAND_31[39:0];
  _RAND_32 = {2{`RANDOM}};
  _T_251 = _RAND_32[39:0];
  _RAND_33 = {2{`RANDOM}};
  _T_254 = _RAND_33[39:0];
  _RAND_34 = {2{`RANDOM}};
  _T_257 = _RAND_34[39:0];
  _RAND_35 = {2{`RANDOM}};
  _T_260 = _RAND_35[39:0];
  _RAND_36 = {2{`RANDOM}};
  _T_263 = _RAND_36[39:0];
  _RAND_37 = {2{`RANDOM}};
  _T_266 = _RAND_37[39:0];
  _RAND_38 = {2{`RANDOM}};
  _T_269 = _RAND_38[39:0];
  _RAND_39 = {2{`RANDOM}};
  _T_272 = _RAND_39[39:0];
  _RAND_40 = {2{`RANDOM}};
  _T_275 = _RAND_40[39:0];
  _RAND_41 = {2{`RANDOM}};
  _T_278 = _RAND_41[39:0];
  _RAND_42 = {2{`RANDOM}};
  _T_281 = _RAND_42[39:0];
  _RAND_43 = {2{`RANDOM}};
  _T_284 = _RAND_43[39:0];
  _RAND_44 = {2{`RANDOM}};
  _T_287 = _RAND_44[39:0];
  _RAND_45 = {2{`RANDOM}};
  _T_290 = _RAND_45[39:0];
  _RAND_46 = {2{`RANDOM}};
  _T_293 = _RAND_46[39:0];
  _RAND_47 = {1{`RANDOM}};
  reg_dpc = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  reg_dscratch = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  reg_dcsr_ebreakm = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  reg_dcsr_step = _RAND_50[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      reg_mstatus_mpie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else if (wen) begin
      if (_T_499) begin
        reg_mstatus_mpie <= _T_1270[7];
      end else begin
        reg_mstatus_mpie <= _GEN_10;
      end
    end else begin
      reg_mstatus_mpie <= _GEN_10;
    end
    if (metaReset) begin
      reg_mstatus_mie <= 1'h0;
    end else if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else if (wen) begin
      if (_T_499) begin
        reg_mstatus_mie <= _T_1270[3];
      end else if (_T_981) begin
        reg_mstatus_mie <= reg_mstatus_mpie;
      end
    end else if (_T_981) begin
      reg_mstatus_mie <= reg_mstatus_mpie;
    end
    if (metaReset) begin
      reg_mepc <= 32'h0;
    end else begin
      reg_mepc <= _GEN_148[31:0];
    end
    if (metaReset) begin
      reg_mcause <= 32'h0;
    end else if (wen) begin
      if (_T_513) begin
        reg_mcause <= _T_1516;
      end else if (insn_break) begin
        reg_mcause <= 32'h3;
      end else if (insn_call) begin
        reg_mcause <= 32'hb;
      end else if (io_exception) begin
        reg_mcause <= 32'h2;
      end
    end else if (insn_break) begin
      reg_mcause <= 32'h3;
    end else if (insn_call) begin
      reg_mcause <= 32'hb;
    end else if (io_exception) begin
      reg_mcause <= 32'h2;
    end
    if (metaReset) begin
      reg_mtval <= 32'h0;
    end else if (wen) begin
      if (_T_511) begin
        reg_mtval <= wdata;
      end
    end
    if (metaReset) begin
      reg_mscratch <= 32'h0;
    end else if (wen) begin
      if (_T_507) begin
        reg_mscratch <= wdata;
      end
    end
    if (metaReset) begin
      reg_medeleg <= 32'h0;
    end else if (wen) begin
      if (_T_523) begin
        reg_medeleg <= wdata;
      end
    end
    if (metaReset) begin
      reg_mip_mtip <= 1'h0;
    end else if (reset) begin
      reg_mip_mtip <= 1'h0;
    end else begin
      reg_mip_mtip <= 1'h1;
    end
    if (metaReset) begin
      reg_mip_msip <= 1'h0;
    end else if (reset) begin
      reg_mip_msip <= 1'h0;
    end else if (wen) begin
      if (_T_503) begin
        reg_mip_msip <= wdata[3];
      end
    end
    if (metaReset) begin
      reg_mie_mtip <= 1'h0;
    end else if (reset) begin
      reg_mie_mtip <= 1'h0;
    end else if (wen) begin
      if (_T_505) begin
        reg_mie_mtip <= wdata[7];
      end
    end
    if (metaReset) begin
      reg_mie_msip <= 1'h0;
    end else if (reset) begin
      reg_mie_msip <= 1'h0;
    end else if (wen) begin
      if (_T_505) begin
        reg_mie_msip <= wdata[3];
      end
    end
    if (metaReset) begin
      _T_176 <= 6'h0;
    end else if (reset) begin
      _T_176 <= 6'h0;
    end else begin
      _T_176 <= _GEN_142[5:0];
    end
    if (metaReset) begin
      _T_180 <= 58'h0;
    end else if (reset) begin
      _T_180 <= 58'h0;
    end else if (wen) begin
      if (_T_487) begin
        _T_180 <= _T_1501[63:6];
      end else if (_T_653) begin
        _T_180 <= _T_1498[63:6];
      end else if (_T_177[6]) begin
        _T_180 <= _T_184;
      end
    end else if (_T_177[6]) begin
      _T_180 <= _T_184;
    end
    if (metaReset) begin
      _T_188 <= 6'h0;
    end else if (reset) begin
      _T_188 <= 6'h0;
    end else begin
      _T_188 <= _GEN_144[5:0];
    end
    if (metaReset) begin
      _T_192 <= 58'h0;
    end else if (reset) begin
      _T_192 <= 58'h0;
    end else if (wen) begin
      if (_T_489) begin
        _T_192 <= _T_1508[63:6];
      end else if (_T_655) begin
        _T_192 <= _T_1505[63:6];
      end else if (_T_189[6]) begin
        _T_192 <= _T_196;
      end
    end else if (_T_189[6]) begin
      _T_192 <= _T_196;
    end
    if (metaReset) begin
      _T_200 <= 40'h0;
    end else begin
      _T_200 <= _GEN_110[39:0];
    end
    if (metaReset) begin
      _T_203 <= 40'h0;
    end else begin
      _T_203 <= _GEN_111[39:0];
    end
    if (metaReset) begin
      _T_206 <= 40'h0;
    end else begin
      _T_206 <= _GEN_112[39:0];
    end
    if (metaReset) begin
      _T_209 <= 40'h0;
    end else begin
      _T_209 <= _GEN_113[39:0];
    end
    if (metaReset) begin
      _T_212 <= 40'h0;
    end else begin
      _T_212 <= _GEN_114[39:0];
    end
    if (metaReset) begin
      _T_215 <= 40'h0;
    end else begin
      _T_215 <= _GEN_115[39:0];
    end
    if (metaReset) begin
      _T_218 <= 40'h0;
    end else begin
      _T_218 <= _GEN_116[39:0];
    end
    if (metaReset) begin
      _T_221 <= 40'h0;
    end else begin
      _T_221 <= _GEN_117[39:0];
    end
    if (metaReset) begin
      _T_224 <= 40'h0;
    end else begin
      _T_224 <= _GEN_118[39:0];
    end
    if (metaReset) begin
      _T_227 <= 40'h0;
    end else begin
      _T_227 <= _GEN_119[39:0];
    end
    if (metaReset) begin
      _T_230 <= 40'h0;
    end else begin
      _T_230 <= _GEN_120[39:0];
    end
    if (metaReset) begin
      _T_233 <= 40'h0;
    end else begin
      _T_233 <= _GEN_121[39:0];
    end
    if (metaReset) begin
      _T_236 <= 40'h0;
    end else begin
      _T_236 <= _GEN_122[39:0];
    end
    if (metaReset) begin
      _T_239 <= 40'h0;
    end else begin
      _T_239 <= _GEN_123[39:0];
    end
    if (metaReset) begin
      _T_242 <= 40'h0;
    end else begin
      _T_242 <= _GEN_124[39:0];
    end
    if (metaReset) begin
      _T_245 <= 40'h0;
    end else begin
      _T_245 <= _GEN_125[39:0];
    end
    if (metaReset) begin
      _T_248 <= 40'h0;
    end else begin
      _T_248 <= _GEN_126[39:0];
    end
    if (metaReset) begin
      _T_251 <= 40'h0;
    end else begin
      _T_251 <= _GEN_127[39:0];
    end
    if (metaReset) begin
      _T_254 <= 40'h0;
    end else begin
      _T_254 <= _GEN_128[39:0];
    end
    if (metaReset) begin
      _T_257 <= 40'h0;
    end else begin
      _T_257 <= _GEN_129[39:0];
    end
    if (metaReset) begin
      _T_260 <= 40'h0;
    end else begin
      _T_260 <= _GEN_130[39:0];
    end
    if (metaReset) begin
      _T_263 <= 40'h0;
    end else begin
      _T_263 <= _GEN_131[39:0];
    end
    if (metaReset) begin
      _T_266 <= 40'h0;
    end else begin
      _T_266 <= _GEN_132[39:0];
    end
    if (metaReset) begin
      _T_269 <= 40'h0;
    end else begin
      _T_269 <= _GEN_133[39:0];
    end
    if (metaReset) begin
      _T_272 <= 40'h0;
    end else begin
      _T_272 <= _GEN_134[39:0];
    end
    if (metaReset) begin
      _T_275 <= 40'h0;
    end else begin
      _T_275 <= _GEN_135[39:0];
    end
    if (metaReset) begin
      _T_278 <= 40'h0;
    end else begin
      _T_278 <= _GEN_136[39:0];
    end
    if (metaReset) begin
      _T_281 <= 40'h0;
    end else begin
      _T_281 <= _GEN_137[39:0];
    end
    if (metaReset) begin
      _T_284 <= 40'h0;
    end else begin
      _T_284 <= _GEN_138[39:0];
    end
    if (metaReset) begin
      _T_287 <= 40'h0;
    end else begin
      _T_287 <= _GEN_139[39:0];
    end
    if (metaReset) begin
      _T_290 <= 40'h0;
    end else begin
      _T_290 <= _GEN_140[39:0];
    end
    if (metaReset) begin
      _T_293 <= 40'h0;
    end else begin
      _T_293 <= _GEN_141[39:0];
    end
    if (metaReset) begin
      reg_dpc <= 32'h0;
    end else if (wen) begin
      if (_T_519) begin
        reg_dpc <= wdata;
      end
    end
    if (metaReset) begin
      reg_dscratch <= 32'h0;
    end else if (wen) begin
      if (_T_521) begin
        reg_dscratch <= wdata;
      end
    end
    if (metaReset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else if (reset) begin
      reg_dcsr_ebreakm <= 1'h0;
    end else if (wen) begin
      if (_T_517) begin
        reg_dcsr_ebreakm <= wdata[15];
      end
    end
    if (metaReset) begin
      reg_dcsr_step <= 1'h0;
    end else if (reset) begin
      reg_dcsr_step <= 1'h0;
    end else if (wen) begin
      if (_T_517) begin
        reg_dcsr_step <= wdata[2];
      end
    end
  end
endmodule
module DatPath(
  input         metaReset,
  input         clock,
  input         reset,
  output [31:0] io_imem_req_bits_pc,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [31:0] io_imem_resp_bits_pc,
  input  [31:0] io_imem_resp_bits_inst,
  output [31:0] io_dmem_req_bits_addr,
  output [31:0] io_dmem_req_bits_data,
  output        io_dmem_req_bits_fcn,
  output [2:0]  io_dmem_req_bits_typ,
  input  [31:0] io_dmem_resp_bits_data,
  input         io_ctl_exe_kill,
  input  [2:0]  io_ctl_pc_sel,
  input         io_ctl_brjmp_sel,
  input  [1:0]  io_ctl_op1_sel,
  input  [1:0]  io_ctl_op2_sel,
  input  [3:0]  io_ctl_alu_fun,
  input  [1:0]  io_ctl_wb_sel,
  input         io_ctl_rf_wen,
  input         io_ctl_bypassable,
  input  [2:0]  io_ctl_csr_cmd,
  input         io_ctl_dmem_fcn,
  input  [2:0]  io_ctl_dmem_typ,
  input         io_ctl_exception,
  output        io_dat_br_eq,
  output        io_dat_br_lt,
  output        io_dat_br_ltu,
  output        io_dat_csr_eret,
  output        _GEN_411,
  output        _GEN_405,
  output        _GEN_426,
  output        _GEN_291,
  output        _GEN_306,
  output        _GEN_384,
  output        _GEN_16_0,
  output        _GEN_19_0,
  output        _GEN_327,
  output        _GEN_390,
  output        _GEN_10_0,
  output        _GEN_285,
  output        _GEN_318,
  output        _GEN_312,
  output        _GEN_399,
  output        _GEN_387,
  output        _GEN_300,
  output        _GEN_279,
  output        _GEN_269,
  output        _GEN_378,
  output        _GEN_368,
  output        _GEN_377,
  output        _GEN_22_0,
  output        _GEN_12_0,
  output        _GEN_294,
  output        _GEN_393,
  output        _GEN_362,
  output        _GEN_461,
  output        _GEN_263,
  output        _GEN_449,
  output        _GEN_288,
  output        _GEN_245,
  output        _GEN_0_0,
  output        _GEN_272,
  output        _GEN_381,
  output        _GEN_371,
  output        _GEN_266,
  output        _GEN_16_1,
  output        _GEN_344,
  output        _GEN_282,
  output        _GEN_443,
  output        _GEN_251,
  output        _GEN_6_0,
  output        _GEN_350,
  output        _GEN_365,
  output        _GEN_15_0,
  output        _GEN_152,
  output        _GEN_446,
  output        _GEN_332,
  output        _GEN_326,
  output        _GEN_359,
  output        _GEN_15_1,
  output        _GEN_458,
  output        _GEN_452,
  output        _GEN_3_0,
  output        _GEN_347,
  output        _GEN_425,
  output        _GEN_239,
  output        _GEN_431,
  output        _GEN_254,
  output        _GEN_353,
  output        _GEN_260,
  output        _GEN_275,
  output        _GEN_9_0,
  output        _GEN_338,
  output        _GEN_374,
  output        _GEN_242,
  output        _GEN_455,
  output        _GEN_413,
  output        _GEN_236,
  output        _GEN_335,
  output        _GEN_18_0,
  output        _GEN_434,
  output        _GEN_248_0,
  output        _GEN_257,
  output        _GEN_320_0,
  output        _GEN_356,
  output        _GEN_12_1,
  output        _GEN_419,
  output        _GEN_314_0,
  output        _GEN_341,
  output        _GEN_440,
  output        _GEN_299_0,
  output        _GEN_398,
  output        _GEN_407,
  output        _GEN_149_0,
  output        _GEN_416,
  output        _GEN_281,
  output        _GEN_15_2,
  output        _GEN_380,
  output        _GEN_296_0,
  output        _GEN_422,
  output        _GEN_329,
  output        _GEN_6_1,
  output        _GEN_437,
  output        _GEN_302_0,
  output        _GEN_401,
  output        _GEN_395,
  output        _GEN_428,
  output        _GEN_308_0,
  output        _GEN_323,
  output        _GEN_317,
  output        _GEN_404,
  output        _GEN_290,
  output        _GEN_9_1,
  output        _GEN_367,
  output        _GEN_284,
  output        _GEN_274_0,
  output        _GEN_383,
  output        _GEN_373,
  output        _GEN_18_2,
  output        _GEN_410,
  output        _GEN_305_0,
  output        _GEN_8_0,
  output        _GEN_2_0,
  output        _GEN_311_0,
  output        _GEN_389,
  output        _GEN_268_0,
  output        _GEN_376,
  output        _GEN_454,
  output        _GEN_293_0,
  output        _GEN_392,
  output        _GEN_361,
  output        _GEN_287,
  output        _GEN_256_0,
  output        _GEN_460,
  output        _GEN_278,
  output        _GEN_355,
  output        _GEN_386,
  output        _GEN_277_0,
  output        _GEN_21_0,
  output        _GEN_262_0,
  output        _GEN_11_0,
  output        _GEN_244_0,
  output        _GEN_448,
  output        _GEN_442,
  output        _GEN_457,
  output        _GEN_337,
  output        _GEN_364,
  output        _GEN_328,
  output        _GEN_463,
  output        _GEN_436,
  output        _GEN_370,
  output        _GEN_250_0,
  output        _GEN_265_0,
  output        _GEN_5_0,
  output        _GEN_271_0,
  output        _GEN_349,
  output        _GEN_343,
  output        _GEN_147,
  output        _GEN_352,
  output        _GEN_247_0,
  output        _GEN_325,
  output        _GEN_151_0,
  output        _GEN_238_0,
  output        _GEN_451,
  output        _GEN_346,
  output        _GEN_409,
  output        _GEN_253_0,
  output        _GEN_331,
  output        _GEN_8_1,
  output        _GEN_11_1,
  output        _GEN_430,
  output        _GEN_424,
  output        _GEN_445,
  output        _GEN_310_0,
  output        _GEN_259_0,
  output        _GEN_358,
  output        _GEN_334,
  output        _GEN_412,
  output        _GEN_11_2,
  output        _GEN_418,
  output        _GEN_427,
  output        _GEN_313_0,
  output        _GEN_292_0,
  output        _GEN_241_0,
  output        _GEN_340,
  output        _GEN_235_0,
  output        _GEN_439,
  output        _GEN_20_0,
  output        _GEN_298_0,
  output        _GEN_307_0,
  output        _GEN_17_0,
  output        _GEN_406,
  output        _GEN_433,
  output        _GEN_319_0,
  output        _GEN_391,
  output        _GEN_400,
  output        _GEN_415,
  output        _GEN_295_0,
  output        _GEN_270_0,
  output        _GEN_4_2,
  output        _GEN_322_0,
  output        _GEN_14_0,
  output        _GEN_421,
  output        _GEN_280_0,
  output        _GEN_379,
  output        _GEN_394,
  output        _GEN_23_0,
  output        _GEN_369,
  output        _GEN_5_2,
  output        _GEN_14_1,
  output        _GEN_13_2,
  output        _GEN_316_0,
  output        _GEN_301_0,
  output        _GEN_283_0,
  output        _GEN_273_0,
  output        _GEN_382,
  output        _GEN_258_0,
  output        _GEN_304_0,
  output        _GEN_403,
  output        _GEN_372,
  output        _GEN_366,
  output        _GEN_267_0,
  output        _GEN_289_0,
  output        _GEN_1_3,
  output        _GEN_388,
  output        _GEN_397,
  output        _GEN_252_0,
  output        _GEN_450,
  output        _GEN_351,
  output        _GEN_17_2,
  output        _GEN_7_2,
  output        _GEN_453,
  output        _GEN_447,
  output        _GEN_438,
  output        _GEN_333,
  output        _GEN_240_0,
  output        _GEN_339,
  output        _GEN_375,
  output        _GEN_261_0,
  output        _GEN_255_0,
  output        _GEN_10_3,
  output        _GEN_360,
  output        _GEN_432,
  output        _GEN_286_0,
  output        _GEN_276_0,
  output        _GEN_459,
  output        _GEN_385,
  output        _GEN_354,
  output        _GEN_234_0,
  output        _GEN_3_3,
  output        _GEN_146,
  output        _GEN_441,
  output        _GEN_321_0,
  output        _GEN_13_3,
  output        _GEN_348,
  output        _GEN_357,
  output        _GEN_243_0,
  output        _GEN_462,
  output        _GEN_456,
  output        _GEN_342,
  output        _GEN_420,
  output        _GEN_414,
  output        _GEN_336,
  output        _GEN_435,
  output        _GEN_249_0,
  output        _GEN_237_0,
  output        _GEN_315_0,
  output        _GEN_264_0,
  output        _GEN_363,
  output        _GEN_246_0,
  output        _GEN_150_0,
  output        _GEN_330,
  output        _GEN_7_3,
  output        _GEN_297_0,
  output        _GEN_345,
  output        _GEN_396,
  output        _GEN_408,
  output        _GEN_423,
  output        _GEN_309_0,
  output        _GEN_303_0,
  output        _GEN_417,
  output        _GEN_429,
  output        _GEN_444,
  output        _GEN_324,
  output        _GEN_402
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire  mem_sparse_metaReset;
  wire  mem_sparse_clock;
  wire  mem_sparse_reset;
  wire [4:0] mem_sparse_io_w_1_addr;
  wire  mem_sparse_io_w_1_en;
  wire [31:0] mem_sparse_io_w_1_data;
  wire [4:0] mem_sparse_io_r_1_addr;
  wire [31:0] mem_sparse_io_r_1_data;
  wire [4:0] mem_sparse_io_r_2_addr;
  wire [31:0] mem_sparse_io_r_2_data;
  wire [3:0] alu_io_fn; // @[dpath.scala 167:20]
  wire [31:0] alu_io_in2; // @[dpath.scala 167:20]
  wire [31:0] alu_io_in1; // @[dpath.scala 167:20]
  wire [31:0] alu_io_out; // @[dpath.scala 167:20]
  wire [31:0] alu_io_adder_out; // @[dpath.scala 167:20]
  wire  alu__GEN_16_0; // @[dpath.scala 167:20]
  wire  alu__GEN_10_0; // @[dpath.scala 167:20]
  wire  alu__GEN_15_1; // @[dpath.scala 167:20]
  wire  alu__GEN_18_0; // @[dpath.scala 167:20]
  wire  alu__GEN_12_1; // @[dpath.scala 167:20]
  wire  alu__GEN_9_1; // @[dpath.scala 167:20]
  wire  alu__GEN_8_1; // @[dpath.scala 167:20]
  wire  alu__GEN_11_2; // @[dpath.scala 167:20]
  wire  alu__GEN_17_0; // @[dpath.scala 167:20]
  wire  alu__GEN_14_0; // @[dpath.scala 167:20]
  wire  alu__GEN_13_3; // @[dpath.scala 167:20]
  wire  csr_metaReset; // @[dpath.scala 216:20]
  wire  csr_clock; // @[dpath.scala 216:20]
  wire  csr_reset; // @[dpath.scala 216:20]
  wire [2:0] csr_io_rw_cmd; // @[dpath.scala 216:20]
  wire [31:0] csr_io_rw_rdata; // @[dpath.scala 216:20]
  wire [31:0] csr_io_rw_wdata; // @[dpath.scala 216:20]
  wire  csr_io_eret; // @[dpath.scala 216:20]
  wire [11:0] csr_io_decode_csr; // @[dpath.scala 216:20]
  wire  csr_io_status_debug; // @[dpath.scala 216:20]
  wire [1:0] csr_io_status_prv; // @[dpath.scala 216:20]
  wire  csr_io_status_sd; // @[dpath.scala 216:20]
  wire [7:0] csr_io_status_zero1; // @[dpath.scala 216:20]
  wire  csr_io_status_tsr; // @[dpath.scala 216:20]
  wire  csr_io_status_tw; // @[dpath.scala 216:20]
  wire  csr_io_status_tvm; // @[dpath.scala 216:20]
  wire  csr_io_status_mxr; // @[dpath.scala 216:20]
  wire  csr_io_status_sum; // @[dpath.scala 216:20]
  wire  csr_io_status_mprv; // @[dpath.scala 216:20]
  wire [1:0] csr_io_status_xs; // @[dpath.scala 216:20]
  wire [1:0] csr_io_status_fs; // @[dpath.scala 216:20]
  wire [1:0] csr_io_status_mpp; // @[dpath.scala 216:20]
  wire [1:0] csr_io_status_hpp; // @[dpath.scala 216:20]
  wire  csr_io_status_spp; // @[dpath.scala 216:20]
  wire  csr_io_status_mpie; // @[dpath.scala 216:20]
  wire  csr_io_status_hpie; // @[dpath.scala 216:20]
  wire  csr_io_status_spie; // @[dpath.scala 216:20]
  wire  csr_io_status_upie; // @[dpath.scala 216:20]
  wire  csr_io_status_mie; // @[dpath.scala 216:20]
  wire  csr_io_status_hie; // @[dpath.scala 216:20]
  wire  csr_io_status_sie; // @[dpath.scala 216:20]
  wire  csr_io_status_uie; // @[dpath.scala 216:20]
  wire [31:0] csr_io_evec; // @[dpath.scala 216:20]
  wire  csr_io_exception; // @[dpath.scala 216:20]
  wire  csr_io_retire; // @[dpath.scala 216:20]
  wire [31:0] csr_io_pc; // @[dpath.scala 216:20]
  wire  csr__GEN_411_0; // @[dpath.scala 216:20]
  wire  csr__GEN_405_0; // @[dpath.scala 216:20]
  wire  csr__GEN_426_0; // @[dpath.scala 216:20]
  wire  csr__GEN_291_0; // @[dpath.scala 216:20]
  wire  csr__GEN_306_0; // @[dpath.scala 216:20]
  wire  csr__GEN_384_0; // @[dpath.scala 216:20]
  wire  csr__GEN_327_0; // @[dpath.scala 216:20]
  wire  csr__GEN_390_0; // @[dpath.scala 216:20]
  wire  csr__GEN_285_0; // @[dpath.scala 216:20]
  wire  csr__GEN_318_0; // @[dpath.scala 216:20]
  wire  csr__GEN_312_0; // @[dpath.scala 216:20]
  wire  csr__GEN_399_0; // @[dpath.scala 216:20]
  wire  csr__GEN_387_0; // @[dpath.scala 216:20]
  wire  csr__GEN_300_0; // @[dpath.scala 216:20]
  wire  csr__GEN_279_0; // @[dpath.scala 216:20]
  wire  csr__GEN_269_0; // @[dpath.scala 216:20]
  wire  csr__GEN_378_0; // @[dpath.scala 216:20]
  wire  csr__GEN_368_0; // @[dpath.scala 216:20]
  wire  csr__GEN_377_0; // @[dpath.scala 216:20]
  wire  csr__GEN_294_0; // @[dpath.scala 216:20]
  wire  csr__GEN_393_0; // @[dpath.scala 216:20]
  wire  csr__GEN_362_0; // @[dpath.scala 216:20]
  wire  csr__GEN_461_0; // @[dpath.scala 216:20]
  wire  csr__GEN_263_0; // @[dpath.scala 216:20]
  wire  csr__GEN_449_0; // @[dpath.scala 216:20]
  wire  csr__GEN_288_0; // @[dpath.scala 216:20]
  wire  csr__GEN_245_0; // @[dpath.scala 216:20]
  wire  csr__GEN_272_0; // @[dpath.scala 216:20]
  wire  csr__GEN_381_0; // @[dpath.scala 216:20]
  wire  csr__GEN_371_0; // @[dpath.scala 216:20]
  wire  csr__GEN_266_0; // @[dpath.scala 216:20]
  wire  csr__GEN_344_0; // @[dpath.scala 216:20]
  wire  csr__GEN_282_0; // @[dpath.scala 216:20]
  wire  csr__GEN_443_0; // @[dpath.scala 216:20]
  wire  csr__GEN_251_0; // @[dpath.scala 216:20]
  wire  csr__GEN_350_0; // @[dpath.scala 216:20]
  wire  csr__GEN_365_0; // @[dpath.scala 216:20]
  wire  csr__GEN_15_0; // @[dpath.scala 216:20]
  wire  csr__GEN_152_0; // @[dpath.scala 216:20]
  wire  csr__GEN_446_0; // @[dpath.scala 216:20]
  wire  csr__GEN_332_0; // @[dpath.scala 216:20]
  wire  csr__GEN_326_0; // @[dpath.scala 216:20]
  wire  csr__GEN_359_0; // @[dpath.scala 216:20]
  wire  csr__GEN_458_0; // @[dpath.scala 216:20]
  wire  csr__GEN_452_0; // @[dpath.scala 216:20]
  wire  csr__GEN_347_0; // @[dpath.scala 216:20]
  wire  csr__GEN_425_0; // @[dpath.scala 216:20]
  wire  csr__GEN_239_0; // @[dpath.scala 216:20]
  wire  csr__GEN_431_0; // @[dpath.scala 216:20]
  wire  csr__GEN_254_0; // @[dpath.scala 216:20]
  wire  csr__GEN_353_0; // @[dpath.scala 216:20]
  wire  csr__GEN_260_0; // @[dpath.scala 216:20]
  wire  csr__GEN_275_0; // @[dpath.scala 216:20]
  wire  csr__GEN_338_0; // @[dpath.scala 216:20]
  wire  csr__GEN_374_0; // @[dpath.scala 216:20]
  wire  csr__GEN_242_0; // @[dpath.scala 216:20]
  wire  csr__GEN_455_0; // @[dpath.scala 216:20]
  wire  csr__GEN_413_0; // @[dpath.scala 216:20]
  wire  csr__GEN_236_0; // @[dpath.scala 216:20]
  wire  csr__GEN_335_0; // @[dpath.scala 216:20]
  wire  csr__GEN_434_0; // @[dpath.scala 216:20]
  wire  csr__GEN_248_1; // @[dpath.scala 216:20]
  wire  csr__GEN_257_0; // @[dpath.scala 216:20]
  wire  csr__GEN_320_1; // @[dpath.scala 216:20]
  wire  csr__GEN_356_0; // @[dpath.scala 216:20]
  wire  csr__GEN_419_0; // @[dpath.scala 216:20]
  wire  csr__GEN_314_1; // @[dpath.scala 216:20]
  wire  csr__GEN_341_0; // @[dpath.scala 216:20]
  wire  csr__GEN_440_0; // @[dpath.scala 216:20]
  wire  csr__GEN_299_1; // @[dpath.scala 216:20]
  wire  csr__GEN_398_0; // @[dpath.scala 216:20]
  wire  csr__GEN_407_0; // @[dpath.scala 216:20]
  wire  csr__GEN_149_1; // @[dpath.scala 216:20]
  wire  csr__GEN_416_0; // @[dpath.scala 216:20]
  wire  csr__GEN_281_0; // @[dpath.scala 216:20]
  wire  csr__GEN_380_0; // @[dpath.scala 216:20]
  wire  csr__GEN_296_1; // @[dpath.scala 216:20]
  wire  csr__GEN_422_0; // @[dpath.scala 216:20]
  wire  csr__GEN_329_0; // @[dpath.scala 216:20]
  wire  csr__GEN_6_1; // @[dpath.scala 216:20]
  wire  csr__GEN_437_0; // @[dpath.scala 216:20]
  wire  csr__GEN_302_1; // @[dpath.scala 216:20]
  wire  csr__GEN_401_0; // @[dpath.scala 216:20]
  wire  csr__GEN_395_0; // @[dpath.scala 216:20]
  wire  csr__GEN_428_0; // @[dpath.scala 216:20]
  wire  csr__GEN_308_1; // @[dpath.scala 216:20]
  wire  csr__GEN_323_0; // @[dpath.scala 216:20]
  wire  csr__GEN_317_0; // @[dpath.scala 216:20]
  wire  csr__GEN_404_0; // @[dpath.scala 216:20]
  wire  csr__GEN_290_0; // @[dpath.scala 216:20]
  wire  csr__GEN_367_0; // @[dpath.scala 216:20]
  wire  csr__GEN_284_0; // @[dpath.scala 216:20]
  wire  csr__GEN_274_1; // @[dpath.scala 216:20]
  wire  csr__GEN_383_0; // @[dpath.scala 216:20]
  wire  csr__GEN_373_0; // @[dpath.scala 216:20]
  wire  csr__GEN_410_0; // @[dpath.scala 216:20]
  wire  csr__GEN_305_1; // @[dpath.scala 216:20]
  wire  csr__GEN_311_1; // @[dpath.scala 216:20]
  wire  csr__GEN_389_0; // @[dpath.scala 216:20]
  wire  csr__GEN_268_1; // @[dpath.scala 216:20]
  wire  csr__GEN_376_0; // @[dpath.scala 216:20]
  wire  csr__GEN_454_0; // @[dpath.scala 216:20]
  wire  csr__GEN_293_1; // @[dpath.scala 216:20]
  wire  csr__GEN_392_0; // @[dpath.scala 216:20]
  wire  csr__GEN_361_0; // @[dpath.scala 216:20]
  wire  csr__GEN_287_0; // @[dpath.scala 216:20]
  wire  csr__GEN_256_1; // @[dpath.scala 216:20]
  wire  csr__GEN_460_0; // @[dpath.scala 216:20]
  wire  csr__GEN_278_0; // @[dpath.scala 216:20]
  wire  csr__GEN_355_0; // @[dpath.scala 216:20]
  wire  csr__GEN_386_0; // @[dpath.scala 216:20]
  wire  csr__GEN_277_1; // @[dpath.scala 216:20]
  wire  csr__GEN_262_1; // @[dpath.scala 216:20]
  wire  csr__GEN_244_1; // @[dpath.scala 216:20]
  wire  csr__GEN_448_0; // @[dpath.scala 216:20]
  wire  csr__GEN_442_0; // @[dpath.scala 216:20]
  wire  csr__GEN_457_0; // @[dpath.scala 216:20]
  wire  csr__GEN_337_0; // @[dpath.scala 216:20]
  wire  csr__GEN_364_0; // @[dpath.scala 216:20]
  wire  csr__GEN_328_0; // @[dpath.scala 216:20]
  wire  csr__GEN_463_0; // @[dpath.scala 216:20]
  wire  csr__GEN_436_0; // @[dpath.scala 216:20]
  wire  csr__GEN_370_0; // @[dpath.scala 216:20]
  wire  csr__GEN_250_1; // @[dpath.scala 216:20]
  wire  csr__GEN_265_1; // @[dpath.scala 216:20]
  wire  csr__GEN_271_1; // @[dpath.scala 216:20]
  wire  csr__GEN_349_0; // @[dpath.scala 216:20]
  wire  csr__GEN_343_0; // @[dpath.scala 216:20]
  wire  csr__GEN_147_0; // @[dpath.scala 216:20]
  wire  csr__GEN_352_0; // @[dpath.scala 216:20]
  wire  csr__GEN_247_1; // @[dpath.scala 216:20]
  wire  csr__GEN_325_0; // @[dpath.scala 216:20]
  wire  csr__GEN_151_1; // @[dpath.scala 216:20]
  wire  csr__GEN_238_1; // @[dpath.scala 216:20]
  wire  csr__GEN_451_0; // @[dpath.scala 216:20]
  wire  csr__GEN_346_0; // @[dpath.scala 216:20]
  wire  csr__GEN_409_0; // @[dpath.scala 216:20]
  wire  csr__GEN_253_1; // @[dpath.scala 216:20]
  wire  csr__GEN_331_0; // @[dpath.scala 216:20]
  wire  csr__GEN_11_1; // @[dpath.scala 216:20]
  wire  csr__GEN_430_0; // @[dpath.scala 216:20]
  wire  csr__GEN_424_0; // @[dpath.scala 216:20]
  wire  csr__GEN_445_0; // @[dpath.scala 216:20]
  wire  csr__GEN_310_1; // @[dpath.scala 216:20]
  wire  csr__GEN_259_1; // @[dpath.scala 216:20]
  wire  csr__GEN_358_0; // @[dpath.scala 216:20]
  wire  csr__GEN_334_0; // @[dpath.scala 216:20]
  wire  csr__GEN_412_0; // @[dpath.scala 216:20]
  wire  csr__GEN_418_0; // @[dpath.scala 216:20]
  wire  csr__GEN_427_0; // @[dpath.scala 216:20]
  wire  csr__GEN_313_1; // @[dpath.scala 216:20]
  wire  csr__GEN_292_1; // @[dpath.scala 216:20]
  wire  csr__GEN_241_1; // @[dpath.scala 216:20]
  wire  csr__GEN_340_0; // @[dpath.scala 216:20]
  wire  csr__GEN_235_1; // @[dpath.scala 216:20]
  wire  csr__GEN_439_0; // @[dpath.scala 216:20]
  wire  csr__GEN_298_1; // @[dpath.scala 216:20]
  wire  csr__GEN_307_1; // @[dpath.scala 216:20]
  wire  csr__GEN_406_0; // @[dpath.scala 216:20]
  wire  csr__GEN_433_0; // @[dpath.scala 216:20]
  wire  csr__GEN_319_1; // @[dpath.scala 216:20]
  wire  csr__GEN_391_0; // @[dpath.scala 216:20]
  wire  csr__GEN_400_0; // @[dpath.scala 216:20]
  wire  csr__GEN_415_0; // @[dpath.scala 216:20]
  wire  csr__GEN_295_1; // @[dpath.scala 216:20]
  wire  csr__GEN_270_1; // @[dpath.scala 216:20]
  wire  csr__GEN_322_1; // @[dpath.scala 216:20]
  wire  csr__GEN_421_0; // @[dpath.scala 216:20]
  wire  csr__GEN_280_1; // @[dpath.scala 216:20]
  wire  csr__GEN_379_0; // @[dpath.scala 216:20]
  wire  csr__GEN_394_0; // @[dpath.scala 216:20]
  wire  csr__GEN_369_0; // @[dpath.scala 216:20]
  wire  csr__GEN_5_2; // @[dpath.scala 216:20]
  wire  csr__GEN_316_1; // @[dpath.scala 216:20]
  wire  csr__GEN_301_1; // @[dpath.scala 216:20]
  wire  csr__GEN_283_1; // @[dpath.scala 216:20]
  wire  csr__GEN_273_1; // @[dpath.scala 216:20]
  wire  csr__GEN_382_0; // @[dpath.scala 216:20]
  wire  csr__GEN_258_1; // @[dpath.scala 216:20]
  wire  csr__GEN_304_1; // @[dpath.scala 216:20]
  wire  csr__GEN_403_0; // @[dpath.scala 216:20]
  wire  csr__GEN_372_0; // @[dpath.scala 216:20]
  wire  csr__GEN_366_0; // @[dpath.scala 216:20]
  wire  csr__GEN_267_1; // @[dpath.scala 216:20]
  wire  csr__GEN_289_1; // @[dpath.scala 216:20]
  wire  csr__GEN_388_0; // @[dpath.scala 216:20]
  wire  csr__GEN_397_0; // @[dpath.scala 216:20]
  wire  csr__GEN_252_1; // @[dpath.scala 216:20]
  wire  csr__GEN_450_0; // @[dpath.scala 216:20]
  wire  csr__GEN_351_0; // @[dpath.scala 216:20]
  wire  csr__GEN_453_0; // @[dpath.scala 216:20]
  wire  csr__GEN_447_0; // @[dpath.scala 216:20]
  wire  csr__GEN_438_0; // @[dpath.scala 216:20]
  wire  csr__GEN_333_0; // @[dpath.scala 216:20]
  wire  csr__GEN_240_1; // @[dpath.scala 216:20]
  wire  csr__GEN_339_0; // @[dpath.scala 216:20]
  wire  csr__GEN_375_0; // @[dpath.scala 216:20]
  wire  csr__GEN_261_1; // @[dpath.scala 216:20]
  wire  csr__GEN_255_1; // @[dpath.scala 216:20]
  wire  csr__GEN_360_0; // @[dpath.scala 216:20]
  wire  csr__GEN_432_0; // @[dpath.scala 216:20]
  wire  csr__GEN_286_1; // @[dpath.scala 216:20]
  wire  csr__GEN_276_1; // @[dpath.scala 216:20]
  wire  csr__GEN_459_0; // @[dpath.scala 216:20]
  wire  csr__GEN_385_0; // @[dpath.scala 216:20]
  wire  csr__GEN_354_0; // @[dpath.scala 216:20]
  wire  csr__GEN_234_1; // @[dpath.scala 216:20]
  wire  csr__GEN_3_3; // @[dpath.scala 216:20]
  wire  csr__GEN_146_0; // @[dpath.scala 216:20]
  wire  csr__GEN_441_0; // @[dpath.scala 216:20]
  wire  csr__GEN_321_1; // @[dpath.scala 216:20]
  wire  csr__GEN_348_0; // @[dpath.scala 216:20]
  wire  csr__GEN_357_0; // @[dpath.scala 216:20]
  wire  csr__GEN_243_1; // @[dpath.scala 216:20]
  wire  csr__GEN_462_0; // @[dpath.scala 216:20]
  wire  csr__GEN_456_0; // @[dpath.scala 216:20]
  wire  csr__GEN_342_0; // @[dpath.scala 216:20]
  wire  csr__GEN_420_0; // @[dpath.scala 216:20]
  wire  csr__GEN_414_0; // @[dpath.scala 216:20]
  wire  csr__GEN_336_0; // @[dpath.scala 216:20]
  wire  csr__GEN_435_0; // @[dpath.scala 216:20]
  wire  csr__GEN_249_1; // @[dpath.scala 216:20]
  wire  csr__GEN_237_1; // @[dpath.scala 216:20]
  wire  csr__GEN_315_1; // @[dpath.scala 216:20]
  wire  csr__GEN_264_1; // @[dpath.scala 216:20]
  wire  csr__GEN_363_0; // @[dpath.scala 216:20]
  wire  csr__GEN_246_1; // @[dpath.scala 216:20]
  wire  csr__GEN_150_1; // @[dpath.scala 216:20]
  wire  csr__GEN_330_0; // @[dpath.scala 216:20]
  wire  csr__GEN_7_3; // @[dpath.scala 216:20]
  wire  csr__GEN_297_1; // @[dpath.scala 216:20]
  wire  csr__GEN_345_0; // @[dpath.scala 216:20]
  wire  csr__GEN_396_0; // @[dpath.scala 216:20]
  wire  csr__GEN_408_0; // @[dpath.scala 216:20]
  wire  csr__GEN_423_0; // @[dpath.scala 216:20]
  wire  csr__GEN_309_1; // @[dpath.scala 216:20]
  wire  csr__GEN_303_1; // @[dpath.scala 216:20]
  wire  csr__GEN_417_0; // @[dpath.scala 216:20]
  wire  csr__GEN_429_0; // @[dpath.scala 216:20]
  wire  csr__GEN_444_0; // @[dpath.scala 216:20]
  wire  csr__GEN_324_0; // @[dpath.scala 216:20]
  wire  csr__GEN_402_0; // @[dpath.scala 216:20]
  reg  wb_reg_valid; // @[dpath.scala 52:29]
  reg [1:0] wb_reg_ctrl_wb_sel; // @[dpath.scala 53:29]
  reg  wb_reg_ctrl_rf_wen; // @[dpath.scala 53:29]
  reg  wb_reg_ctrl_bypassable; // @[dpath.scala 53:29]
  reg [2:0] wb_reg_ctrl_csr_cmd; // @[dpath.scala 53:29]
  reg [31:0] wb_reg_alu; // @[dpath.scala 54:29]
  reg [11:0] wb_reg_csr_addr; // @[dpath.scala 55:29]
  reg [4:0] wb_reg_wbaddr; // @[dpath.scala 56:29]
  wire [4:0] exe_rs1_addr = io_imem_resp_bits_inst[19:15]; // @[dpath.scala 83:31]
  wire  _T_129 = wb_reg_wbaddr == exe_rs1_addr; // @[dpath.scala 105:42]
  wire  _T_131 = exe_rs1_addr != 5'h0; // @[dpath.scala 105:77]
  wire  _T_132 = _T_129 & _T_131; // @[dpath.scala 105:60]
  wire  _T_133 = _T_132 & wb_reg_ctrl_rf_wen; // @[dpath.scala 105:85]
  wire  _T_135 = ~wb_reg_ctrl_bypassable; // @[dpath.scala 105:110]
  wire  _T_136 = _T_133 & _T_135; // @[dpath.scala 105:107]
  wire [4:0] exe_rs2_addr = io_imem_resp_bits_inst[24:20]; // @[dpath.scala 84:31]
  wire  _T_137 = wb_reg_wbaddr == exe_rs2_addr; // @[dpath.scala 106:42]
  wire  _T_139 = exe_rs2_addr != 5'h0; // @[dpath.scala 106:77]
  wire  _T_140 = _T_137 & _T_139; // @[dpath.scala 106:60]
  wire  _T_141 = _T_140 & wb_reg_ctrl_rf_wen; // @[dpath.scala 106:85]
  wire  _T_144 = _T_141 & _T_135; // @[dpath.scala 106:107]
  wire  wb_hazard_stall = _T_136 | _T_144; // @[dpath.scala 105:135]
  wire  _T_124 = ~wb_hazard_stall; // @[dpath.scala 66:26]
  wire  _T_125 = io_ctl_pc_sel == 3'h4; // @[dpath.scala 69:36]
  wire  _T_126 = io_ctl_pc_sel == 3'h3; // @[dpath.scala 70:36]
  wire [31:0] exe_jump_reg_target = alu_io_adder_out; // @[dpath.scala 63:34 dpath.scala 178:24]
  wire [19:0] imm_j = {io_imem_resp_bits_inst[31],io_imem_resp_bits_inst[19:12],io_imem_resp_bits_inst[20],io_imem_resp_bits_inst[30:21]}; // @[Cat.scala 30:58]
  wire [10:0] _T_203 = imm_j[19] ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12]
  wire [31:0] imm_j_sext = {_T_203,io_imem_resp_bits_inst[31],io_imem_resp_bits_inst[19:12],io_imem_resp_bits_inst[20],io_imem_resp_bits_inst[30:21],1'h0}; // @[Cat.scala 30:58]
  wire [11:0] imm_b = {io_imem_resp_bits_inst[31],io_imem_resp_bits_inst[7],io_imem_resp_bits_inst[30:25],io_imem_resp_bits_inst[11:8]}; // @[Cat.scala 30:58]
  wire [18:0] _T_196 = imm_b[11] ? 19'h7ffff : 19'h0; // @[Bitwise.scala 72:12]
  wire [31:0] imm_b_sext = {_T_196,io_imem_resp_bits_inst[31],io_imem_resp_bits_inst[7],io_imem_resp_bits_inst[30:25],io_imem_resp_bits_inst[11:8],1'h0}; // @[Cat.scala 30:58]
  wire [31:0] imm_brjmp = io_ctl_brjmp_sel ? imm_j_sext : imm_b_sext; // @[dpath.scala 176:23]
  wire [31:0] exe_brjmp_target = io_imem_resp_bits_pc + imm_brjmp; // @[dpath.scala 177:31]
  wire [31:0] _T_127 = _T_126 ? exe_jump_reg_target : exe_brjmp_target; // @[dpath.scala 70:21]
  wire [31:0] exception_target = csr_io_evec; // @[dpath.scala 64:34 dpath.scala 226:21]
  wire [4:0] exe_wbaddr = io_imem_resp_bits_inst[11:7]; // @[dpath.scala 85:31]
  wire  _T_151 = wb_reg_wbaddr != 5'h0; // @[dpath.scala 121:47]
  wire  _T_311 = wb_reg_ctrl_wb_sel == 2'h0; // @[dpath.scala 238:39]
  wire  _T_312 = wb_reg_ctrl_wb_sel == 2'h1; // @[dpath.scala 239:39]
  wire  _T_313 = wb_reg_ctrl_wb_sel == 2'h2; // @[dpath.scala 240:39]
  wire  _T_314 = wb_reg_ctrl_wb_sel == 2'h3; // @[dpath.scala 241:39]
  wire [31:0] _T_315 = _T_314 ? csr_io_rw_rdata : wb_reg_alu; // @[Mux.scala 61:16]
  wire [31:0] _T_316 = _T_313 ? io_imem_resp_bits_pc : _T_315; // @[Mux.scala 61:16]
  wire [31:0] _T_317 = _T_312 ? io_dmem_resp_bits_data : _T_316; // @[Mux.scala 61:16]
  wire [31:0] regfile__T_156_data = mem_sparse_io_r_1_data;
  wire [31:0] rf_rs1_data = _T_131 ? regfile__T_156_data : 32'h0; // @[dpath.scala 126:25]
  wire [31:0] regfile__T_160_data = mem_sparse_io_r_2_data;
  wire [31:0] rf_rs2_data = _T_139 ? regfile__T_160_data : 32'h0; // @[dpath.scala 127:25]
  wire [11:0] imm_i = io_imem_resp_bits_inst[31:20]; // @[dpath.scala 131:24]
  wire [11:0] imm_s = {io_imem_resp_bits_inst[31:25],exe_wbaddr}; // @[Cat.scala 30:58]
  wire [31:0] imm_u = {io_imem_resp_bits_inst[31:12],12'h0}; // @[Cat.scala 30:58]
  wire [19:0] _T_186 = imm_i[11] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [31:0] imm_i_sext = {_T_186,imm_i}; // @[Cat.scala 30:58]
  wire [19:0] _T_191 = imm_s[11] ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12]
  wire [31:0] imm_s_sext = {_T_191,io_imem_resp_bits_inst[31:25],exe_wbaddr}; // @[Cat.scala 30:58]
  wire  _T_211 = _T_133 & wb_reg_ctrl_bypassable; // @[dpath.scala 148:109]
  wire [31:0] exe_rs1_data = _T_211 ? wb_reg_alu : rf_rs1_data; // @[Mux.scala 61:16]
  wire  _T_217 = _T_141 & wb_reg_ctrl_bypassable; // @[dpath.scala 151:109]
  wire [31:0] exe_rs2_data = _T_217 ? wb_reg_alu : rf_rs2_data; // @[Mux.scala 61:16]
  wire  _T_218 = io_ctl_op1_sel == 2'h2; // @[dpath.scala 156:41]
  wire  _T_219 = io_ctl_op1_sel == 2'h1; // @[dpath.scala 157:41]
  wire [31:0] _T_220 = _T_219 ? imm_u : exe_rs1_data; // @[dpath.scala 157:25]
  wire  _T_221 = io_ctl_op2_sel == 2'h1; // @[dpath.scala 160:41]
  wire  _T_222 = io_ctl_op2_sel == 2'h3; // @[dpath.scala 161:41]
  wire  _T_223 = io_ctl_op2_sel == 2'h2; // @[dpath.scala 162:41]
  wire [31:0] _T_224 = _T_223 ? imm_s_sext : exe_rs2_data; // @[dpath.scala 162:25]
  wire [31:0] _T_225 = _T_222 ? io_imem_resp_bits_pc : _T_224; // @[dpath.scala 161:25]
  wire [31:0] _T_229 = _T_211 ? wb_reg_alu : rf_rs1_data;
  wire [31:0] _T_230 = _T_217 ? wb_reg_alu : rf_rs2_data;
  wire  _T_235 = io_ctl_dmem_fcn & _T_124; // @[dpath.scala 191:48]
  wire  _T_237 = wb_hazard_stall | io_ctl_exe_kill; // @[dpath.scala 199:26]
  wire  _T_244 = io_imem_resp_valid & _T_124; // @[dpath.scala 213:30]
  reg  _T_246; // @[dpath.scala 224:27]
  SparseMem mem_sparse (
    .metaReset(mem_sparse_metaReset),
    .clock(mem_sparse_clock),
    .reset(mem_sparse_reset),
    .io_w_1_addr(mem_sparse_io_w_1_addr),
    .io_w_1_en(mem_sparse_io_w_1_en),
    .io_w_1_data(mem_sparse_io_w_1_data),
    .io_r_1_addr(mem_sparse_io_r_1_addr),
    .io_r_1_data(mem_sparse_io_r_1_data),
    .io_r_2_addr(mem_sparse_io_r_2_addr),
    .io_r_2_data(mem_sparse_io_r_2_data)
  );
  ALU alu ( // @[dpath.scala 167:20]
    .io_fn(alu_io_fn),
    .io_in2(alu_io_in2),
    .io_in1(alu_io_in1),
    .io_out(alu_io_out),
    .io_adder_out(alu_io_adder_out),
    ._GEN_16_0(alu__GEN_16_0),
    ._GEN_10_0(alu__GEN_10_0),
    ._GEN_15_1(alu__GEN_15_1),
    ._GEN_18_0(alu__GEN_18_0),
    ._GEN_12_1(alu__GEN_12_1),
    ._GEN_9_1(alu__GEN_9_1),
    ._GEN_8_1(alu__GEN_8_1),
    ._GEN_11_2(alu__GEN_11_2),
    ._GEN_17_0(alu__GEN_17_0),
    ._GEN_14_0(alu__GEN_14_0),
    ._GEN_13_3(alu__GEN_13_3)
  );
  CSRFile csr ( // @[dpath.scala 216:20]
    .metaReset(csr_metaReset),
    .clock(csr_clock),
    .reset(csr_reset),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_eret(csr_io_eret),
    .io_decode_csr(csr_io_decode_csr),
    .io_status_debug(csr_io_status_debug),
    .io_status_prv(csr_io_status_prv),
    .io_status_sd(csr_io_status_sd),
    .io_status_zero1(csr_io_status_zero1),
    .io_status_tsr(csr_io_status_tsr),
    .io_status_tw(csr_io_status_tw),
    .io_status_tvm(csr_io_status_tvm),
    .io_status_mxr(csr_io_status_mxr),
    .io_status_sum(csr_io_status_sum),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_xs(csr_io_status_xs),
    .io_status_fs(csr_io_status_fs),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_hpp(csr_io_status_hpp),
    .io_status_spp(csr_io_status_spp),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_hpie(csr_io_status_hpie),
    .io_status_spie(csr_io_status_spie),
    .io_status_upie(csr_io_status_upie),
    .io_status_mie(csr_io_status_mie),
    .io_status_hie(csr_io_status_hie),
    .io_status_sie(csr_io_status_sie),
    .io_status_uie(csr_io_status_uie),
    .io_evec(csr_io_evec),
    .io_exception(csr_io_exception),
    .io_retire(csr_io_retire),
    .io_pc(csr_io_pc),
    ._GEN_411_0(csr__GEN_411_0),
    ._GEN_405_0(csr__GEN_405_0),
    ._GEN_426_0(csr__GEN_426_0),
    ._GEN_291_0(csr__GEN_291_0),
    ._GEN_306_0(csr__GEN_306_0),
    ._GEN_384_0(csr__GEN_384_0),
    ._GEN_327_0(csr__GEN_327_0),
    ._GEN_390_0(csr__GEN_390_0),
    ._GEN_285_0(csr__GEN_285_0),
    ._GEN_318_0(csr__GEN_318_0),
    ._GEN_312_0(csr__GEN_312_0),
    ._GEN_399_0(csr__GEN_399_0),
    ._GEN_387_0(csr__GEN_387_0),
    ._GEN_300_0(csr__GEN_300_0),
    ._GEN_279_0(csr__GEN_279_0),
    ._GEN_269_0(csr__GEN_269_0),
    ._GEN_378_0(csr__GEN_378_0),
    ._GEN_368_0(csr__GEN_368_0),
    ._GEN_377_0(csr__GEN_377_0),
    ._GEN_294_0(csr__GEN_294_0),
    ._GEN_393_0(csr__GEN_393_0),
    ._GEN_362_0(csr__GEN_362_0),
    ._GEN_461_0(csr__GEN_461_0),
    ._GEN_263_0(csr__GEN_263_0),
    ._GEN_449_0(csr__GEN_449_0),
    ._GEN_288_0(csr__GEN_288_0),
    ._GEN_245_0(csr__GEN_245_0),
    ._GEN_272_0(csr__GEN_272_0),
    ._GEN_381_0(csr__GEN_381_0),
    ._GEN_371_0(csr__GEN_371_0),
    ._GEN_266_0(csr__GEN_266_0),
    ._GEN_344_0(csr__GEN_344_0),
    ._GEN_282_0(csr__GEN_282_0),
    ._GEN_443_0(csr__GEN_443_0),
    ._GEN_251_0(csr__GEN_251_0),
    ._GEN_350_0(csr__GEN_350_0),
    ._GEN_365_0(csr__GEN_365_0),
    ._GEN_15_0(csr__GEN_15_0),
    ._GEN_152_0(csr__GEN_152_0),
    ._GEN_446_0(csr__GEN_446_0),
    ._GEN_332_0(csr__GEN_332_0),
    ._GEN_326_0(csr__GEN_326_0),
    ._GEN_359_0(csr__GEN_359_0),
    ._GEN_458_0(csr__GEN_458_0),
    ._GEN_452_0(csr__GEN_452_0),
    ._GEN_347_0(csr__GEN_347_0),
    ._GEN_425_0(csr__GEN_425_0),
    ._GEN_239_0(csr__GEN_239_0),
    ._GEN_431_0(csr__GEN_431_0),
    ._GEN_254_0(csr__GEN_254_0),
    ._GEN_353_0(csr__GEN_353_0),
    ._GEN_260_0(csr__GEN_260_0),
    ._GEN_275_0(csr__GEN_275_0),
    ._GEN_338_0(csr__GEN_338_0),
    ._GEN_374_0(csr__GEN_374_0),
    ._GEN_242_0(csr__GEN_242_0),
    ._GEN_455_0(csr__GEN_455_0),
    ._GEN_413_0(csr__GEN_413_0),
    ._GEN_236_0(csr__GEN_236_0),
    ._GEN_335_0(csr__GEN_335_0),
    ._GEN_434_0(csr__GEN_434_0),
    ._GEN_248_1(csr__GEN_248_1),
    ._GEN_257_0(csr__GEN_257_0),
    ._GEN_320_1(csr__GEN_320_1),
    ._GEN_356_0(csr__GEN_356_0),
    ._GEN_419_0(csr__GEN_419_0),
    ._GEN_314_1(csr__GEN_314_1),
    ._GEN_341_0(csr__GEN_341_0),
    ._GEN_440_0(csr__GEN_440_0),
    ._GEN_299_1(csr__GEN_299_1),
    ._GEN_398_0(csr__GEN_398_0),
    ._GEN_407_0(csr__GEN_407_0),
    ._GEN_149_1(csr__GEN_149_1),
    ._GEN_416_0(csr__GEN_416_0),
    ._GEN_281_0(csr__GEN_281_0),
    ._GEN_380_0(csr__GEN_380_0),
    ._GEN_296_1(csr__GEN_296_1),
    ._GEN_422_0(csr__GEN_422_0),
    ._GEN_329_0(csr__GEN_329_0),
    ._GEN_6_1(csr__GEN_6_1),
    ._GEN_437_0(csr__GEN_437_0),
    ._GEN_302_1(csr__GEN_302_1),
    ._GEN_401_0(csr__GEN_401_0),
    ._GEN_395_0(csr__GEN_395_0),
    ._GEN_428_0(csr__GEN_428_0),
    ._GEN_308_1(csr__GEN_308_1),
    ._GEN_323_0(csr__GEN_323_0),
    ._GEN_317_0(csr__GEN_317_0),
    ._GEN_404_0(csr__GEN_404_0),
    ._GEN_290_0(csr__GEN_290_0),
    ._GEN_367_0(csr__GEN_367_0),
    ._GEN_284_0(csr__GEN_284_0),
    ._GEN_274_1(csr__GEN_274_1),
    ._GEN_383_0(csr__GEN_383_0),
    ._GEN_373_0(csr__GEN_373_0),
    ._GEN_410_0(csr__GEN_410_0),
    ._GEN_305_1(csr__GEN_305_1),
    ._GEN_311_1(csr__GEN_311_1),
    ._GEN_389_0(csr__GEN_389_0),
    ._GEN_268_1(csr__GEN_268_1),
    ._GEN_376_0(csr__GEN_376_0),
    ._GEN_454_0(csr__GEN_454_0),
    ._GEN_293_1(csr__GEN_293_1),
    ._GEN_392_0(csr__GEN_392_0),
    ._GEN_361_0(csr__GEN_361_0),
    ._GEN_287_0(csr__GEN_287_0),
    ._GEN_256_1(csr__GEN_256_1),
    ._GEN_460_0(csr__GEN_460_0),
    ._GEN_278_0(csr__GEN_278_0),
    ._GEN_355_0(csr__GEN_355_0),
    ._GEN_386_0(csr__GEN_386_0),
    ._GEN_277_1(csr__GEN_277_1),
    ._GEN_262_1(csr__GEN_262_1),
    ._GEN_244_1(csr__GEN_244_1),
    ._GEN_448_0(csr__GEN_448_0),
    ._GEN_442_0(csr__GEN_442_0),
    ._GEN_457_0(csr__GEN_457_0),
    ._GEN_337_0(csr__GEN_337_0),
    ._GEN_364_0(csr__GEN_364_0),
    ._GEN_328_0(csr__GEN_328_0),
    ._GEN_463_0(csr__GEN_463_0),
    ._GEN_436_0(csr__GEN_436_0),
    ._GEN_370_0(csr__GEN_370_0),
    ._GEN_250_1(csr__GEN_250_1),
    ._GEN_265_1(csr__GEN_265_1),
    ._GEN_271_1(csr__GEN_271_1),
    ._GEN_349_0(csr__GEN_349_0),
    ._GEN_343_0(csr__GEN_343_0),
    ._GEN_147_0(csr__GEN_147_0),
    ._GEN_352_0(csr__GEN_352_0),
    ._GEN_247_1(csr__GEN_247_1),
    ._GEN_325_0(csr__GEN_325_0),
    ._GEN_151_1(csr__GEN_151_1),
    ._GEN_238_1(csr__GEN_238_1),
    ._GEN_451_0(csr__GEN_451_0),
    ._GEN_346_0(csr__GEN_346_0),
    ._GEN_409_0(csr__GEN_409_0),
    ._GEN_253_1(csr__GEN_253_1),
    ._GEN_331_0(csr__GEN_331_0),
    ._GEN_11_1(csr__GEN_11_1),
    ._GEN_430_0(csr__GEN_430_0),
    ._GEN_424_0(csr__GEN_424_0),
    ._GEN_445_0(csr__GEN_445_0),
    ._GEN_310_1(csr__GEN_310_1),
    ._GEN_259_1(csr__GEN_259_1),
    ._GEN_358_0(csr__GEN_358_0),
    ._GEN_334_0(csr__GEN_334_0),
    ._GEN_412_0(csr__GEN_412_0),
    ._GEN_418_0(csr__GEN_418_0),
    ._GEN_427_0(csr__GEN_427_0),
    ._GEN_313_1(csr__GEN_313_1),
    ._GEN_292_1(csr__GEN_292_1),
    ._GEN_241_1(csr__GEN_241_1),
    ._GEN_340_0(csr__GEN_340_0),
    ._GEN_235_1(csr__GEN_235_1),
    ._GEN_439_0(csr__GEN_439_0),
    ._GEN_298_1(csr__GEN_298_1),
    ._GEN_307_1(csr__GEN_307_1),
    ._GEN_406_0(csr__GEN_406_0),
    ._GEN_433_0(csr__GEN_433_0),
    ._GEN_319_1(csr__GEN_319_1),
    ._GEN_391_0(csr__GEN_391_0),
    ._GEN_400_0(csr__GEN_400_0),
    ._GEN_415_0(csr__GEN_415_0),
    ._GEN_295_1(csr__GEN_295_1),
    ._GEN_270_1(csr__GEN_270_1),
    ._GEN_322_1(csr__GEN_322_1),
    ._GEN_421_0(csr__GEN_421_0),
    ._GEN_280_1(csr__GEN_280_1),
    ._GEN_379_0(csr__GEN_379_0),
    ._GEN_394_0(csr__GEN_394_0),
    ._GEN_369_0(csr__GEN_369_0),
    ._GEN_5_2(csr__GEN_5_2),
    ._GEN_316_1(csr__GEN_316_1),
    ._GEN_301_1(csr__GEN_301_1),
    ._GEN_283_1(csr__GEN_283_1),
    ._GEN_273_1(csr__GEN_273_1),
    ._GEN_382_0(csr__GEN_382_0),
    ._GEN_258_1(csr__GEN_258_1),
    ._GEN_304_1(csr__GEN_304_1),
    ._GEN_403_0(csr__GEN_403_0),
    ._GEN_372_0(csr__GEN_372_0),
    ._GEN_366_0(csr__GEN_366_0),
    ._GEN_267_1(csr__GEN_267_1),
    ._GEN_289_1(csr__GEN_289_1),
    ._GEN_388_0(csr__GEN_388_0),
    ._GEN_397_0(csr__GEN_397_0),
    ._GEN_252_1(csr__GEN_252_1),
    ._GEN_450_0(csr__GEN_450_0),
    ._GEN_351_0(csr__GEN_351_0),
    ._GEN_453_0(csr__GEN_453_0),
    ._GEN_447_0(csr__GEN_447_0),
    ._GEN_438_0(csr__GEN_438_0),
    ._GEN_333_0(csr__GEN_333_0),
    ._GEN_240_1(csr__GEN_240_1),
    ._GEN_339_0(csr__GEN_339_0),
    ._GEN_375_0(csr__GEN_375_0),
    ._GEN_261_1(csr__GEN_261_1),
    ._GEN_255_1(csr__GEN_255_1),
    ._GEN_360_0(csr__GEN_360_0),
    ._GEN_432_0(csr__GEN_432_0),
    ._GEN_286_1(csr__GEN_286_1),
    ._GEN_276_1(csr__GEN_276_1),
    ._GEN_459_0(csr__GEN_459_0),
    ._GEN_385_0(csr__GEN_385_0),
    ._GEN_354_0(csr__GEN_354_0),
    ._GEN_234_1(csr__GEN_234_1),
    ._GEN_3_3(csr__GEN_3_3),
    ._GEN_146_0(csr__GEN_146_0),
    ._GEN_441_0(csr__GEN_441_0),
    ._GEN_321_1(csr__GEN_321_1),
    ._GEN_348_0(csr__GEN_348_0),
    ._GEN_357_0(csr__GEN_357_0),
    ._GEN_243_1(csr__GEN_243_1),
    ._GEN_462_0(csr__GEN_462_0),
    ._GEN_456_0(csr__GEN_456_0),
    ._GEN_342_0(csr__GEN_342_0),
    ._GEN_420_0(csr__GEN_420_0),
    ._GEN_414_0(csr__GEN_414_0),
    ._GEN_336_0(csr__GEN_336_0),
    ._GEN_435_0(csr__GEN_435_0),
    ._GEN_249_1(csr__GEN_249_1),
    ._GEN_237_1(csr__GEN_237_1),
    ._GEN_315_1(csr__GEN_315_1),
    ._GEN_264_1(csr__GEN_264_1),
    ._GEN_363_0(csr__GEN_363_0),
    ._GEN_246_1(csr__GEN_246_1),
    ._GEN_150_1(csr__GEN_150_1),
    ._GEN_330_0(csr__GEN_330_0),
    ._GEN_7_3(csr__GEN_7_3),
    ._GEN_297_1(csr__GEN_297_1),
    ._GEN_345_0(csr__GEN_345_0),
    ._GEN_396_0(csr__GEN_396_0),
    ._GEN_408_0(csr__GEN_408_0),
    ._GEN_423_0(csr__GEN_423_0),
    ._GEN_309_1(csr__GEN_309_1),
    ._GEN_303_1(csr__GEN_303_1),
    ._GEN_417_0(csr__GEN_417_0),
    ._GEN_429_0(csr__GEN_429_0),
    ._GEN_444_0(csr__GEN_444_0),
    ._GEN_324_0(csr__GEN_324_0),
    ._GEN_402_0(csr__GEN_402_0)
  );
  assign mem_sparse_metaReset = metaReset;
  assign csr_metaReset = metaReset;
  assign io_imem_req_bits_pc = _T_125 ? exception_target : _T_127; // @[dpath.scala 73:24]
  assign io_imem_resp_ready = ~wb_hazard_stall; // @[dpath.scala 66:23]
  assign io_dmem_req_bits_addr = alu_io_out; // @[dpath.scala 193:26]
  assign io_dmem_req_bits_data = _T_217 ? wb_reg_alu : rf_rs2_data; // @[dpath.scala 194:26]
  assign io_dmem_req_bits_fcn = _T_235 & io_imem_resp_valid; // @[dpath.scala 191:29]
  assign io_dmem_req_bits_typ = io_ctl_dmem_typ; // @[dpath.scala 192:26]
  assign io_dat_br_eq = exe_rs1_data == exe_rs2_data; // @[dpath.scala 182:18]
  assign io_dat_br_lt = $signed(_T_229) < $signed(_T_230); // @[dpath.scala 183:18]
  assign io_dat_br_ltu = exe_rs1_data < exe_rs2_data; // @[dpath.scala 184:18]
  assign io_dat_csr_eret = csr_io_eret; // @[dpath.scala 227:20]
  assign _GEN_411 = csr__GEN_411_0;
  assign _GEN_405 = csr__GEN_405_0;
  assign _GEN_426 = csr__GEN_426_0;
  assign _GEN_291 = csr__GEN_291_0;
  assign _GEN_306 = csr__GEN_306_0;
  assign _GEN_384 = csr__GEN_384_0;
  assign _GEN_16_0 = alu__GEN_16_0;
  assign _GEN_19_0 = io_ctl_op2_sel == 2'h1;
  assign _GEN_327 = csr__GEN_327_0;
  assign _GEN_390 = csr__GEN_390_0;
  assign _GEN_10_0 = alu__GEN_10_0;
  assign _GEN_285 = csr__GEN_285_0;
  assign _GEN_318 = csr__GEN_318_0;
  assign _GEN_312 = csr__GEN_312_0;
  assign _GEN_399 = csr__GEN_399_0;
  assign _GEN_387 = csr__GEN_387_0;
  assign _GEN_300 = csr__GEN_300_0;
  assign _GEN_279 = csr__GEN_279_0;
  assign _GEN_269 = csr__GEN_269_0;
  assign _GEN_378 = csr__GEN_378_0;
  assign _GEN_368 = csr__GEN_368_0;
  assign _GEN_377 = csr__GEN_377_0;
  assign _GEN_22_0 = wb_hazard_stall | io_ctl_exe_kill;
  assign _GEN_12_0 = _T_141 & wb_reg_ctrl_bypassable;
  assign _GEN_294 = csr__GEN_294_0;
  assign _GEN_393 = csr__GEN_393_0;
  assign _GEN_362 = csr__GEN_362_0;
  assign _GEN_461 = csr__GEN_461_0;
  assign _GEN_263 = csr__GEN_263_0;
  assign _GEN_449 = csr__GEN_449_0;
  assign _GEN_288 = csr__GEN_288_0;
  assign _GEN_245 = csr__GEN_245_0;
  assign _GEN_0_0 = imm_j[19];
  assign _GEN_272 = csr__GEN_272_0;
  assign _GEN_381 = csr__GEN_381_0;
  assign _GEN_371 = csr__GEN_371_0;
  assign _GEN_266 = csr__GEN_266_0;
  assign _GEN_16_1 = io_ctl_pc_sel == 3'h4;
  assign _GEN_344 = csr__GEN_344_0;
  assign _GEN_282 = csr__GEN_282_0;
  assign _GEN_443 = csr__GEN_443_0;
  assign _GEN_251 = csr__GEN_251_0;
  assign _GEN_6_0 = wb_reg_ctrl_wb_sel == 2'h1;
  assign _GEN_350 = csr__GEN_350_0;
  assign _GEN_365 = csr__GEN_365_0;
  assign _GEN_15_0 = csr__GEN_15_0;
  assign _GEN_152 = csr__GEN_152_0;
  assign _GEN_446 = csr__GEN_446_0;
  assign _GEN_332 = csr__GEN_332_0;
  assign _GEN_326 = csr__GEN_326_0;
  assign _GEN_359 = csr__GEN_359_0;
  assign _GEN_15_1 = alu__GEN_15_1;
  assign _GEN_458 = csr__GEN_458_0;
  assign _GEN_452 = csr__GEN_452_0;
  assign _GEN_3_0 = io_ctl_pc_sel == 3'h3;
  assign _GEN_347 = csr__GEN_347_0;
  assign _GEN_425 = csr__GEN_425_0;
  assign _GEN_239 = csr__GEN_239_0;
  assign _GEN_431 = csr__GEN_431_0;
  assign _GEN_254 = csr__GEN_254_0;
  assign _GEN_353 = csr__GEN_353_0;
  assign _GEN_260 = csr__GEN_260_0;
  assign _GEN_275 = csr__GEN_275_0;
  assign _GEN_9_0 = imm_i[11];
  assign _GEN_338 = csr__GEN_338_0;
  assign _GEN_374 = csr__GEN_374_0;
  assign _GEN_242 = csr__GEN_242_0;
  assign _GEN_455 = csr__GEN_455_0;
  assign _GEN_413 = csr__GEN_413_0;
  assign _GEN_236 = csr__GEN_236_0;
  assign _GEN_335 = csr__GEN_335_0;
  assign _GEN_18_0 = alu__GEN_18_0;
  assign _GEN_434 = csr__GEN_434_0;
  assign _GEN_248_0 = csr__GEN_248_1;
  assign _GEN_257 = csr__GEN_257_0;
  assign _GEN_320_0 = csr__GEN_320_1;
  assign _GEN_356 = csr__GEN_356_0;
  assign _GEN_12_1 = alu__GEN_12_1;
  assign _GEN_419 = csr__GEN_419_0;
  assign _GEN_314_0 = csr__GEN_314_1;
  assign _GEN_341 = csr__GEN_341_0;
  assign _GEN_440 = csr__GEN_440_0;
  assign _GEN_299_0 = csr__GEN_299_1;
  assign _GEN_398 = csr__GEN_398_0;
  assign _GEN_407 = csr__GEN_407_0;
  assign _GEN_149_0 = csr__GEN_149_1;
  assign _GEN_416 = csr__GEN_416_0;
  assign _GEN_281 = csr__GEN_281_0;
  assign _GEN_15_2 = io_ctl_op2_sel == 2'h3;
  assign _GEN_380 = csr__GEN_380_0;
  assign _GEN_296_0 = csr__GEN_296_1;
  assign _GEN_422 = csr__GEN_422_0;
  assign _GEN_329 = csr__GEN_329_0;
  assign _GEN_6_1 = csr__GEN_6_1;
  assign _GEN_437 = csr__GEN_437_0;
  assign _GEN_302_0 = csr__GEN_302_1;
  assign _GEN_401 = csr__GEN_401_0;
  assign _GEN_395 = csr__GEN_395_0;
  assign _GEN_428 = csr__GEN_428_0;
  assign _GEN_308_0 = csr__GEN_308_1;
  assign _GEN_323 = csr__GEN_323_0;
  assign _GEN_317 = csr__GEN_317_0;
  assign _GEN_404 = csr__GEN_404_0;
  assign _GEN_290 = csr__GEN_290_0;
  assign _GEN_9_1 = alu__GEN_9_1;
  assign _GEN_367 = csr__GEN_367_0;
  assign _GEN_284 = csr__GEN_284_0;
  assign _GEN_274_0 = csr__GEN_274_1;
  assign _GEN_383 = csr__GEN_383_0;
  assign _GEN_373 = csr__GEN_373_0;
  assign _GEN_18_2 = wb_reg_ctrl_wb_sel == 2'h0;
  assign _GEN_410 = csr__GEN_410_0;
  assign _GEN_305_0 = csr__GEN_305_1;
  assign _GEN_8_0 = exe_rs2_addr != 5'h0;
  assign _GEN_2_0 = io_ctl_brjmp_sel;
  assign _GEN_311_0 = csr__GEN_311_1;
  assign _GEN_389 = csr__GEN_389_0;
  assign _GEN_268_0 = csr__GEN_268_1;
  assign _GEN_376 = csr__GEN_376_0;
  assign _GEN_454 = csr__GEN_454_0;
  assign _GEN_293_0 = csr__GEN_293_1;
  assign _GEN_392 = csr__GEN_392_0;
  assign _GEN_361 = csr__GEN_361_0;
  assign _GEN_287 = csr__GEN_287_0;
  assign _GEN_256_0 = csr__GEN_256_1;
  assign _GEN_460 = csr__GEN_460_0;
  assign _GEN_278 = csr__GEN_278_0;
  assign _GEN_355 = csr__GEN_355_0;
  assign _GEN_386 = csr__GEN_386_0;
  assign _GEN_277_0 = csr__GEN_277_1;
  assign _GEN_21_0 = reset;
  assign _GEN_262_0 = csr__GEN_262_1;
  assign _GEN_11_0 = _T_133 & wb_reg_ctrl_bypassable;
  assign _GEN_244_0 = csr__GEN_244_1;
  assign _GEN_448 = csr__GEN_448_0;
  assign _GEN_442 = csr__GEN_442_0;
  assign _GEN_457 = csr__GEN_457_0;
  assign _GEN_337 = csr__GEN_337_0;
  assign _GEN_364 = csr__GEN_364_0;
  assign _GEN_328 = csr__GEN_328_0;
  assign _GEN_463 = csr__GEN_463_0;
  assign _GEN_436 = csr__GEN_436_0;
  assign _GEN_370 = csr__GEN_370_0;
  assign _GEN_250_0 = csr__GEN_250_1;
  assign _GEN_265_0 = csr__GEN_265_1;
  assign _GEN_5_0 = wb_reg_ctrl_wb_sel == 2'h2;
  assign _GEN_271_0 = csr__GEN_271_1;
  assign _GEN_349 = csr__GEN_349_0;
  assign _GEN_343 = csr__GEN_343_0;
  assign _GEN_147 = csr__GEN_147_0;
  assign _GEN_352 = csr__GEN_352_0;
  assign _GEN_247_0 = csr__GEN_247_1;
  assign _GEN_325 = csr__GEN_325_0;
  assign _GEN_151_0 = csr__GEN_151_1;
  assign _GEN_238_0 = csr__GEN_238_1;
  assign _GEN_451 = csr__GEN_451_0;
  assign _GEN_346 = csr__GEN_346_0;
  assign _GEN_409 = csr__GEN_409_0;
  assign _GEN_253_0 = csr__GEN_253_1;
  assign _GEN_331 = csr__GEN_331_0;
  assign _GEN_8_1 = alu__GEN_8_1;
  assign _GEN_11_1 = csr__GEN_11_1;
  assign _GEN_430 = csr__GEN_430_0;
  assign _GEN_424 = csr__GEN_424_0;
  assign _GEN_445 = csr__GEN_445_0;
  assign _GEN_310_0 = csr__GEN_310_1;
  assign _GEN_259_0 = csr__GEN_259_1;
  assign _GEN_358 = csr__GEN_358_0;
  assign _GEN_334 = csr__GEN_334_0;
  assign _GEN_412 = csr__GEN_412_0;
  assign _GEN_11_2 = alu__GEN_11_2;
  assign _GEN_418 = csr__GEN_418_0;
  assign _GEN_427 = csr__GEN_427_0;
  assign _GEN_313_0 = csr__GEN_313_1;
  assign _GEN_292_0 = csr__GEN_292_1;
  assign _GEN_241_0 = csr__GEN_241_1;
  assign _GEN_340 = csr__GEN_340_0;
  assign _GEN_235_0 = csr__GEN_235_1;
  assign _GEN_439 = csr__GEN_439_0;
  assign _GEN_20_0 = io_ctl_op1_sel == 2'h2;
  assign _GEN_298_0 = csr__GEN_298_1;
  assign _GEN_307_0 = csr__GEN_307_1;
  assign _GEN_17_0 = alu__GEN_17_0;
  assign _GEN_406 = csr__GEN_406_0;
  assign _GEN_433 = csr__GEN_433_0;
  assign _GEN_319_0 = csr__GEN_319_1;
  assign _GEN_391 = csr__GEN_391_0;
  assign _GEN_400 = csr__GEN_400_0;
  assign _GEN_415 = csr__GEN_415_0;
  assign _GEN_295_0 = csr__GEN_295_1;
  assign _GEN_270_0 = csr__GEN_270_1;
  assign _GEN_4_2 = wb_reg_ctrl_wb_sel == 2'h3;
  assign _GEN_322_0 = csr__GEN_322_1;
  assign _GEN_14_0 = alu__GEN_14_0;
  assign _GEN_421 = csr__GEN_421_0;
  assign _GEN_280_0 = csr__GEN_280_1;
  assign _GEN_379 = csr__GEN_379_0;
  assign _GEN_394 = csr__GEN_394_0;
  assign _GEN_23_0 = wb_hazard_stall | io_ctl_exe_kill;
  assign _GEN_369 = csr__GEN_369_0;
  assign _GEN_5_2 = csr__GEN_5_2;
  assign _GEN_14_1 = io_ctl_op2_sel == 2'h2;
  assign _GEN_13_2 = io_ctl_op1_sel == 2'h1;
  assign _GEN_316_0 = csr__GEN_316_1;
  assign _GEN_301_0 = csr__GEN_301_1;
  assign _GEN_283_0 = csr__GEN_283_1;
  assign _GEN_273_0 = csr__GEN_273_1;
  assign _GEN_382 = csr__GEN_382_0;
  assign _GEN_258_0 = csr__GEN_258_1;
  assign _GEN_304_0 = csr__GEN_304_1;
  assign _GEN_403 = csr__GEN_403_0;
  assign _GEN_372 = csr__GEN_372_0;
  assign _GEN_366 = csr__GEN_366_0;
  assign _GEN_267_0 = csr__GEN_267_1;
  assign _GEN_289_0 = csr__GEN_289_1;
  assign _GEN_1_3 = imm_b[11];
  assign _GEN_388 = csr__GEN_388_0;
  assign _GEN_397 = csr__GEN_397_0;
  assign _GEN_252_0 = csr__GEN_252_1;
  assign _GEN_450 = csr__GEN_450_0;
  assign _GEN_351 = csr__GEN_351_0;
  assign _GEN_17_2 = _T_141 & wb_reg_ctrl_bypassable;
  assign _GEN_7_2 = exe_rs1_addr != 5'h0;
  assign _GEN_453 = csr__GEN_453_0;
  assign _GEN_447 = csr__GEN_447_0;
  assign _GEN_438 = csr__GEN_438_0;
  assign _GEN_333 = csr__GEN_333_0;
  assign _GEN_240_0 = csr__GEN_240_1;
  assign _GEN_339 = csr__GEN_339_0;
  assign _GEN_375 = csr__GEN_375_0;
  assign _GEN_261_0 = csr__GEN_261_1;
  assign _GEN_255_0 = csr__GEN_255_1;
  assign _GEN_10_3 = imm_s[11];
  assign _GEN_360 = csr__GEN_360_0;
  assign _GEN_432 = csr__GEN_432_0;
  assign _GEN_286_0 = csr__GEN_286_1;
  assign _GEN_276_0 = csr__GEN_276_1;
  assign _GEN_459 = csr__GEN_459_0;
  assign _GEN_385 = csr__GEN_385_0;
  assign _GEN_354 = csr__GEN_354_0;
  assign _GEN_234_0 = csr__GEN_234_1;
  assign _GEN_3_3 = csr__GEN_3_3;
  assign _GEN_146 = csr__GEN_146_0;
  assign _GEN_441 = csr__GEN_441_0;
  assign _GEN_321_0 = csr__GEN_321_1;
  assign _GEN_13_3 = alu__GEN_13_3;
  assign _GEN_348 = csr__GEN_348_0;
  assign _GEN_357 = csr__GEN_357_0;
  assign _GEN_243_0 = csr__GEN_243_1;
  assign _GEN_462 = csr__GEN_462_0;
  assign _GEN_456 = csr__GEN_456_0;
  assign _GEN_342 = csr__GEN_342_0;
  assign _GEN_420 = csr__GEN_420_0;
  assign _GEN_414 = csr__GEN_414_0;
  assign _GEN_336 = csr__GEN_336_0;
  assign _GEN_435 = csr__GEN_435_0;
  assign _GEN_249_0 = csr__GEN_249_1;
  assign _GEN_237_0 = csr__GEN_237_1;
  assign _GEN_315_0 = csr__GEN_315_1;
  assign _GEN_264_0 = csr__GEN_264_1;
  assign _GEN_363 = csr__GEN_363_0;
  assign _GEN_246_0 = csr__GEN_246_1;
  assign _GEN_150_0 = csr__GEN_150_1;
  assign _GEN_330 = csr__GEN_330_0;
  assign _GEN_7_3 = csr__GEN_7_3;
  assign _GEN_297_0 = csr__GEN_297_1;
  assign _GEN_345 = csr__GEN_345_0;
  assign _GEN_396 = csr__GEN_396_0;
  assign _GEN_408 = csr__GEN_408_0;
  assign _GEN_423 = csr__GEN_423_0;
  assign _GEN_309_0 = csr__GEN_309_1;
  assign _GEN_303_0 = csr__GEN_303_1;
  assign _GEN_417 = csr__GEN_417_0;
  assign _GEN_429 = csr__GEN_429_0;
  assign _GEN_444 = csr__GEN_444_0;
  assign _GEN_324 = csr__GEN_324_0;
  assign _GEN_402 = csr__GEN_402_0;
  assign mem_sparse_clock = clock;
  assign mem_sparse_reset = reset;
  assign mem_sparse_io_w_1_addr = wb_reg_wbaddr;
  assign mem_sparse_io_w_1_en = wb_reg_ctrl_rf_wen & _T_151;
  assign mem_sparse_io_w_1_data = _T_311 ? wb_reg_alu : _T_317;
  assign mem_sparse_io_r_1_addr = io_imem_resp_bits_inst[19:15];
  assign mem_sparse_io_r_2_addr = io_imem_resp_bits_inst[24:20];
  assign alu_io_fn = io_ctl_alu_fun; // @[dpath.scala 171:18]
  assign alu_io_in2 = _T_221 ? imm_i_sext : _T_225; // @[dpath.scala 170:18]
  assign alu_io_in1 = _T_218 ? {{27'd0}, exe_rs1_addr} : _T_220; // @[dpath.scala 169:18]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_rw_cmd = wb_reg_ctrl_csr_cmd; // @[dpath.scala 220:21]
  assign csr_io_rw_wdata = wb_reg_alu; // @[dpath.scala 219:21]
  assign csr_io_decode_csr = wb_reg_csr_addr; // @[dpath.scala 218:24]
  assign csr_io_exception = _T_246; // @[dpath.scala 224:21]
  assign csr_io_retire = wb_reg_valid; // @[dpath.scala 223:21]
  assign csr_io_pc = io_imem_resp_bits_pc - 32'h4; // @[dpath.scala 225:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wb_reg_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wb_reg_ctrl_wb_sel = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  wb_reg_ctrl_rf_wen = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  wb_reg_ctrl_bypassable = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  wb_reg_ctrl_csr_cmd = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  wb_reg_alu = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  wb_reg_csr_addr = _RAND_6[11:0];
  _RAND_7 = {1{`RANDOM}};
  wb_reg_wbaddr = _RAND_7[4:0];
  _RAND_8 = {1{`RANDOM}};
  _T_246 = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      wb_reg_valid <= 1'h0;
    end else if (reset) begin
      wb_reg_valid <= 1'h0;
    end else begin
      wb_reg_valid <= _T_244;
    end
    if (metaReset) begin
      wb_reg_ctrl_wb_sel <= 2'h0;
    end else begin
      wb_reg_ctrl_wb_sel <= io_ctl_wb_sel;
    end
    if (metaReset) begin
      wb_reg_ctrl_rf_wen <= 1'h0;
    end else if (_T_237) begin
      wb_reg_ctrl_rf_wen <= 1'h0;
    end else begin
      wb_reg_ctrl_rf_wen <= io_ctl_rf_wen;
    end
    if (metaReset) begin
      wb_reg_ctrl_bypassable <= 1'h0;
    end else begin
      wb_reg_ctrl_bypassable <= io_ctl_bypassable;
    end
    if (metaReset) begin
      wb_reg_ctrl_csr_cmd <= 3'h0;
    end else if (_T_237) begin
      wb_reg_ctrl_csr_cmd <= 3'h0;
    end else begin
      wb_reg_ctrl_csr_cmd <= io_ctl_csr_cmd;
    end
    if (metaReset) begin
      wb_reg_alu <= 32'h0;
    end else begin
      wb_reg_alu <= alu_io_out;
    end
    if (metaReset) begin
      wb_reg_csr_addr <= 12'h0;
    end else begin
      wb_reg_csr_addr <= io_imem_resp_bits_inst[31:20];
    end
    if (metaReset) begin
      wb_reg_wbaddr <= 5'h0;
    end else begin
      wb_reg_wbaddr <= io_imem_resp_bits_inst[11:7];
    end
    if (metaReset) begin
      _T_246 <= 1'h0;
    end else begin
      _T_246 <= io_ctl_exception;
    end
  end
endmodule
module SparseMem(
  input         metaReset,
  input         clock,
  input         reset,
  input  [4:0]  io_w_1_addr,
  input         io_w_1_en,
  input  [31:0] io_w_1_data,
  input  [4:0]  io_r_1_addr,
  output [31:0] io_r_1_data,
  input  [4:0]  io_r_2_addr,
  output [31:0] io_r_2_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem [0:31];
  wire [31:0] mem__T_152_data;
  wire [4:0] mem__T_152_addr;
  wire [31:0] mem__T_274_data;
  wire [4:0] mem__T_274_addr;
  wire [31:0] mem__T_396_data;
  wire [4:0] mem__T_396_addr;
  wire [31:0] mem__T_528_data;
  wire [4:0] mem__T_528_addr;
  wire  mem__T_528_mask;
  wire  mem__T_528_en;
  wire [31:0] mem__T_656_data;
  wire [4:0] mem__T_656_addr;
  wire  mem__T_656_mask;
  wire  mem__T_656_en;
  reg  addresses_0_valid;
  reg [4:0] addresses_0_bits;
  reg  addresses_1_valid;
  reg [4:0] addresses_1_bits;
  reg  addresses_2_valid;
  reg [4:0] addresses_2_bits;
  reg  addresses_3_valid;
  reg [4:0] addresses_3_bits;
  reg  addresses_4_valid;
  reg [4:0] addresses_4_bits;
  reg  addresses_5_valid;
  reg [4:0] addresses_5_bits;
  reg  addresses_6_valid;
  reg [4:0] addresses_6_bits;
  reg  addresses_7_valid;
  reg [4:0] addresses_7_bits;
  reg  addresses_8_valid;
  reg [4:0] addresses_8_bits;
  reg  addresses_9_valid;
  reg [4:0] addresses_9_bits;
  reg  addresses_10_valid;
  reg [4:0] addresses_10_bits;
  reg  addresses_11_valid;
  reg [4:0] addresses_11_bits;
  reg  addresses_12_valid;
  reg [4:0] addresses_12_bits;
  reg  addresses_13_valid;
  reg [4:0] addresses_13_bits;
  reg  addresses_14_valid;
  reg [4:0] addresses_14_bits;
  reg  addresses_15_valid;
  reg [4:0] addresses_15_bits;
  reg  addresses_16_valid;
  reg [4:0] addresses_16_bits;
  reg  addresses_17_valid;
  reg [4:0] addresses_17_bits;
  reg  addresses_18_valid;
  reg [4:0] addresses_18_bits;
  reg  addresses_19_valid;
  reg [4:0] addresses_19_bits;
  reg  addresses_20_valid;
  reg [4:0] addresses_20_bits;
  reg  addresses_21_valid;
  reg [4:0] addresses_21_bits;
  reg  addresses_22_valid;
  reg [4:0] addresses_22_bits;
  reg  addresses_23_valid;
  reg [4:0] addresses_23_bits;
  reg  addresses_24_valid;
  reg [4:0] addresses_24_bits;
  reg  addresses_25_valid;
  reg [4:0] addresses_25_bits;
  reg  addresses_26_valid;
  reg [4:0] addresses_26_bits;
  reg  addresses_27_valid;
  reg [4:0] addresses_27_bits;
  reg  addresses_28_valid;
  reg [4:0] addresses_28_bits;
  reg  addresses_29_valid;
  reg [4:0] addresses_29_bits;
  reg  addresses_30_valid;
  reg [4:0] addresses_30_bits;
  reg  addresses_31_valid;
  reg [4:0] addresses_31_bits;
  wire  _T_33 = addresses_0_bits == 5'h0;
  wire  _T_34 = addresses_0_valid & _T_33;
  wire  _T_35 = addresses_1_bits == 5'h0;
  wire  _T_36 = addresses_1_valid & _T_35;
  wire  _T_37 = addresses_2_bits == 5'h0;
  wire  _T_38 = addresses_2_valid & _T_37;
  wire  _T_39 = addresses_3_bits == 5'h0;
  wire  _T_40 = addresses_3_valid & _T_39;
  wire  _T_41 = addresses_4_bits == 5'h0;
  wire  _T_42 = addresses_4_valid & _T_41;
  wire  _T_43 = addresses_5_bits == 5'h0;
  wire  _T_44 = addresses_5_valid & _T_43;
  wire  _T_45 = addresses_6_bits == 5'h0;
  wire  _T_46 = addresses_6_valid & _T_45;
  wire  _T_47 = addresses_7_bits == 5'h0;
  wire  _T_48 = addresses_7_valid & _T_47;
  wire  _T_49 = addresses_8_bits == 5'h0;
  wire  _T_50 = addresses_8_valid & _T_49;
  wire  _T_51 = addresses_9_bits == 5'h0;
  wire  _T_52 = addresses_9_valid & _T_51;
  wire  _T_53 = addresses_10_bits == 5'h0;
  wire  _T_54 = addresses_10_valid & _T_53;
  wire  _T_55 = addresses_11_bits == 5'h0;
  wire  _T_56 = addresses_11_valid & _T_55;
  wire  _T_57 = addresses_12_bits == 5'h0;
  wire  _T_58 = addresses_12_valid & _T_57;
  wire  _T_59 = addresses_13_bits == 5'h0;
  wire  _T_60 = addresses_13_valid & _T_59;
  wire  _T_61 = addresses_14_bits == 5'h0;
  wire  _T_62 = addresses_14_valid & _T_61;
  wire  _T_63 = addresses_15_bits == 5'h0;
  wire  _T_64 = addresses_15_valid & _T_63;
  wire  _T_65 = addresses_16_bits == 5'h0;
  wire  _T_66 = addresses_16_valid & _T_65;
  wire  _T_67 = addresses_17_bits == 5'h0;
  wire  _T_68 = addresses_17_valid & _T_67;
  wire  _T_69 = addresses_18_bits == 5'h0;
  wire  _T_70 = addresses_18_valid & _T_69;
  wire  _T_71 = addresses_19_bits == 5'h0;
  wire  _T_72 = addresses_19_valid & _T_71;
  wire  _T_73 = addresses_20_bits == 5'h0;
  wire  _T_74 = addresses_20_valid & _T_73;
  wire  _T_75 = addresses_21_bits == 5'h0;
  wire  _T_76 = addresses_21_valid & _T_75;
  wire  _T_77 = addresses_22_bits == 5'h0;
  wire  _T_78 = addresses_22_valid & _T_77;
  wire  _T_79 = addresses_23_bits == 5'h0;
  wire  _T_80 = addresses_23_valid & _T_79;
  wire  _T_81 = addresses_24_bits == 5'h0;
  wire  _T_82 = addresses_24_valid & _T_81;
  wire  _T_83 = addresses_25_bits == 5'h0;
  wire  _T_84 = addresses_25_valid & _T_83;
  wire  _T_85 = addresses_26_bits == 5'h0;
  wire  _T_86 = addresses_26_valid & _T_85;
  wire  _T_87 = addresses_27_bits == 5'h0;
  wire  _T_88 = addresses_27_valid & _T_87;
  wire  _T_89 = addresses_28_bits == 5'h0;
  wire  _T_90 = addresses_28_valid & _T_89;
  wire  _T_91 = addresses_29_bits == 5'h0;
  wire  _T_92 = addresses_29_valid & _T_91;
  wire  _T_93 = addresses_30_bits == 5'h0;
  wire  _T_94 = addresses_30_valid & _T_93;
  wire  _T_95 = addresses_31_bits == 5'h0;
  wire  _T_96 = addresses_31_valid & _T_95;
  wire [7:0] _T_104 = {_T_48,_T_46,_T_44,_T_42,_T_40,_T_38,_T_36,_T_34};
  wire [15:0] _T_112 = {_T_64,_T_62,_T_60,_T_58,_T_56,_T_54,_T_52,_T_50,_T_104};
  wire [7:0] _T_119 = {_T_80,_T_78,_T_76,_T_74,_T_72,_T_70,_T_68,_T_66};
  wire [31:0] _T_128 = {_T_96,_T_94,_T_92,_T_90,_T_88,_T_86,_T_84,_T_82,_T_119,_T_112};
  wire  _T_129 = _T_128 != 32'h0;
  wire  _T_132 = |_T_128[31:16];
  wire [15:0] _T_133 = _T_128[31:16] | _T_128[15:0];
  wire  _T_136 = |_T_133[15:8];
  wire [7:0] _T_137 = _T_133[15:8] | _T_133[7:0];
  wire  _T_140 = |_T_137[7:4];
  wire [3:0] _T_141 = _T_137[7:4] | _T_137[3:0];
  wire  _T_144 = |_T_141[3:2];
  wire [1:0] _T_145 = _T_141[3:2] | _T_141[1:0];
  wire [3:0] _T_149 = {_T_136,_T_140,_T_144,_T_145[1]};
  wire [4:0] _T_150 = {_T_132,_T_136,_T_140,_T_144,_T_145[1]};
  wire  _T_155 = addresses_0_bits == io_r_1_addr;
  wire  _T_156 = addresses_0_valid & _T_155;
  wire  _T_157 = addresses_1_bits == io_r_1_addr;
  wire  _T_158 = addresses_1_valid & _T_157;
  wire  _T_159 = addresses_2_bits == io_r_1_addr;
  wire  _T_160 = addresses_2_valid & _T_159;
  wire  _T_161 = addresses_3_bits == io_r_1_addr;
  wire  _T_162 = addresses_3_valid & _T_161;
  wire  _T_163 = addresses_4_bits == io_r_1_addr;
  wire  _T_164 = addresses_4_valid & _T_163;
  wire  _T_165 = addresses_5_bits == io_r_1_addr;
  wire  _T_166 = addresses_5_valid & _T_165;
  wire  _T_167 = addresses_6_bits == io_r_1_addr;
  wire  _T_168 = addresses_6_valid & _T_167;
  wire  _T_169 = addresses_7_bits == io_r_1_addr;
  wire  _T_170 = addresses_7_valid & _T_169;
  wire  _T_171 = addresses_8_bits == io_r_1_addr;
  wire  _T_172 = addresses_8_valid & _T_171;
  wire  _T_173 = addresses_9_bits == io_r_1_addr;
  wire  _T_174 = addresses_9_valid & _T_173;
  wire  _T_175 = addresses_10_bits == io_r_1_addr;
  wire  _T_176 = addresses_10_valid & _T_175;
  wire  _T_177 = addresses_11_bits == io_r_1_addr;
  wire  _T_178 = addresses_11_valid & _T_177;
  wire  _T_179 = addresses_12_bits == io_r_1_addr;
  wire  _T_180 = addresses_12_valid & _T_179;
  wire  _T_181 = addresses_13_bits == io_r_1_addr;
  wire  _T_182 = addresses_13_valid & _T_181;
  wire  _T_183 = addresses_14_bits == io_r_1_addr;
  wire  _T_184 = addresses_14_valid & _T_183;
  wire  _T_185 = addresses_15_bits == io_r_1_addr;
  wire  _T_186 = addresses_15_valid & _T_185;
  wire  _T_187 = addresses_16_bits == io_r_1_addr;
  wire  _T_188 = addresses_16_valid & _T_187;
  wire  _T_189 = addresses_17_bits == io_r_1_addr;
  wire  _T_190 = addresses_17_valid & _T_189;
  wire  _T_191 = addresses_18_bits == io_r_1_addr;
  wire  _T_192 = addresses_18_valid & _T_191;
  wire  _T_193 = addresses_19_bits == io_r_1_addr;
  wire  _T_194 = addresses_19_valid & _T_193;
  wire  _T_195 = addresses_20_bits == io_r_1_addr;
  wire  _T_196 = addresses_20_valid & _T_195;
  wire  _T_197 = addresses_21_bits == io_r_1_addr;
  wire  _T_198 = addresses_21_valid & _T_197;
  wire  _T_199 = addresses_22_bits == io_r_1_addr;
  wire  _T_200 = addresses_22_valid & _T_199;
  wire  _T_201 = addresses_23_bits == io_r_1_addr;
  wire  _T_202 = addresses_23_valid & _T_201;
  wire  _T_203 = addresses_24_bits == io_r_1_addr;
  wire  _T_204 = addresses_24_valid & _T_203;
  wire  _T_205 = addresses_25_bits == io_r_1_addr;
  wire  _T_206 = addresses_25_valid & _T_205;
  wire  _T_207 = addresses_26_bits == io_r_1_addr;
  wire  _T_208 = addresses_26_valid & _T_207;
  wire  _T_209 = addresses_27_bits == io_r_1_addr;
  wire  _T_210 = addresses_27_valid & _T_209;
  wire  _T_211 = addresses_28_bits == io_r_1_addr;
  wire  _T_212 = addresses_28_valid & _T_211;
  wire  _T_213 = addresses_29_bits == io_r_1_addr;
  wire  _T_214 = addresses_29_valid & _T_213;
  wire  _T_215 = addresses_30_bits == io_r_1_addr;
  wire  _T_216 = addresses_30_valid & _T_215;
  wire  _T_217 = addresses_31_bits == io_r_1_addr;
  wire  _T_218 = addresses_31_valid & _T_217;
  wire [7:0] _T_226 = {_T_170,_T_168,_T_166,_T_164,_T_162,_T_160,_T_158,_T_156};
  wire [15:0] _T_234 = {_T_186,_T_184,_T_182,_T_180,_T_178,_T_176,_T_174,_T_172,_T_226};
  wire [7:0] _T_241 = {_T_202,_T_200,_T_198,_T_196,_T_194,_T_192,_T_190,_T_188};
  wire [31:0] _T_250 = {_T_218,_T_216,_T_214,_T_212,_T_210,_T_208,_T_206,_T_204,_T_241,_T_234};
  wire  _T_251 = _T_250 != 32'h0;
  wire  _T_254 = |_T_250[31:16];
  wire [15:0] _T_255 = _T_250[31:16] | _T_250[15:0];
  wire  _T_258 = |_T_255[15:8];
  wire [7:0] _T_259 = _T_255[15:8] | _T_255[7:0];
  wire  _T_262 = |_T_259[7:4];
  wire [3:0] _T_263 = _T_259[7:4] | _T_259[3:0];
  wire  _T_266 = |_T_263[3:2];
  wire [1:0] _T_267 = _T_263[3:2] | _T_263[1:0];
  wire [3:0] _T_271 = {_T_258,_T_262,_T_266,_T_267[1]};
  wire  _T_277 = addresses_0_bits == io_r_2_addr;
  wire  _T_278 = addresses_0_valid & _T_277;
  wire  _T_279 = addresses_1_bits == io_r_2_addr;
  wire  _T_280 = addresses_1_valid & _T_279;
  wire  _T_281 = addresses_2_bits == io_r_2_addr;
  wire  _T_282 = addresses_2_valid & _T_281;
  wire  _T_283 = addresses_3_bits == io_r_2_addr;
  wire  _T_284 = addresses_3_valid & _T_283;
  wire  _T_285 = addresses_4_bits == io_r_2_addr;
  wire  _T_286 = addresses_4_valid & _T_285;
  wire  _T_287 = addresses_5_bits == io_r_2_addr;
  wire  _T_288 = addresses_5_valid & _T_287;
  wire  _T_289 = addresses_6_bits == io_r_2_addr;
  wire  _T_290 = addresses_6_valid & _T_289;
  wire  _T_291 = addresses_7_bits == io_r_2_addr;
  wire  _T_292 = addresses_7_valid & _T_291;
  wire  _T_293 = addresses_8_bits == io_r_2_addr;
  wire  _T_294 = addresses_8_valid & _T_293;
  wire  _T_295 = addresses_9_bits == io_r_2_addr;
  wire  _T_296 = addresses_9_valid & _T_295;
  wire  _T_297 = addresses_10_bits == io_r_2_addr;
  wire  _T_298 = addresses_10_valid & _T_297;
  wire  _T_299 = addresses_11_bits == io_r_2_addr;
  wire  _T_300 = addresses_11_valid & _T_299;
  wire  _T_301 = addresses_12_bits == io_r_2_addr;
  wire  _T_302 = addresses_12_valid & _T_301;
  wire  _T_303 = addresses_13_bits == io_r_2_addr;
  wire  _T_304 = addresses_13_valid & _T_303;
  wire  _T_305 = addresses_14_bits == io_r_2_addr;
  wire  _T_306 = addresses_14_valid & _T_305;
  wire  _T_307 = addresses_15_bits == io_r_2_addr;
  wire  _T_308 = addresses_15_valid & _T_307;
  wire  _T_309 = addresses_16_bits == io_r_2_addr;
  wire  _T_310 = addresses_16_valid & _T_309;
  wire  _T_311 = addresses_17_bits == io_r_2_addr;
  wire  _T_312 = addresses_17_valid & _T_311;
  wire  _T_313 = addresses_18_bits == io_r_2_addr;
  wire  _T_314 = addresses_18_valid & _T_313;
  wire  _T_315 = addresses_19_bits == io_r_2_addr;
  wire  _T_316 = addresses_19_valid & _T_315;
  wire  _T_317 = addresses_20_bits == io_r_2_addr;
  wire  _T_318 = addresses_20_valid & _T_317;
  wire  _T_319 = addresses_21_bits == io_r_2_addr;
  wire  _T_320 = addresses_21_valid & _T_319;
  wire  _T_321 = addresses_22_bits == io_r_2_addr;
  wire  _T_322 = addresses_22_valid & _T_321;
  wire  _T_323 = addresses_23_bits == io_r_2_addr;
  wire  _T_324 = addresses_23_valid & _T_323;
  wire  _T_325 = addresses_24_bits == io_r_2_addr;
  wire  _T_326 = addresses_24_valid & _T_325;
  wire  _T_327 = addresses_25_bits == io_r_2_addr;
  wire  _T_328 = addresses_25_valid & _T_327;
  wire  _T_329 = addresses_26_bits == io_r_2_addr;
  wire  _T_330 = addresses_26_valid & _T_329;
  wire  _T_331 = addresses_27_bits == io_r_2_addr;
  wire  _T_332 = addresses_27_valid & _T_331;
  wire  _T_333 = addresses_28_bits == io_r_2_addr;
  wire  _T_334 = addresses_28_valid & _T_333;
  wire  _T_335 = addresses_29_bits == io_r_2_addr;
  wire  _T_336 = addresses_29_valid & _T_335;
  wire  _T_337 = addresses_30_bits == io_r_2_addr;
  wire  _T_338 = addresses_30_valid & _T_337;
  wire  _T_339 = addresses_31_bits == io_r_2_addr;
  wire  _T_340 = addresses_31_valid & _T_339;
  wire [7:0] _T_348 = {_T_292,_T_290,_T_288,_T_286,_T_284,_T_282,_T_280,_T_278};
  wire [15:0] _T_356 = {_T_308,_T_306,_T_304,_T_302,_T_300,_T_298,_T_296,_T_294,_T_348};
  wire [7:0] _T_363 = {_T_324,_T_322,_T_320,_T_318,_T_316,_T_314,_T_312,_T_310};
  wire [31:0] _T_372 = {_T_340,_T_338,_T_336,_T_334,_T_332,_T_330,_T_328,_T_326,_T_363,_T_356};
  wire  _T_373 = _T_372 != 32'h0;
  wire  _T_376 = |_T_372[31:16];
  wire [15:0] _T_377 = _T_372[31:16] | _T_372[15:0];
  wire  _T_380 = |_T_377[15:8];
  wire [7:0] _T_381 = _T_377[15:8] | _T_377[7:0];
  wire  _T_384 = |_T_381[7:4];
  wire [3:0] _T_385 = _T_381[7:4] | _T_381[3:0];
  wire  _T_388 = |_T_385[3:2];
  wire [1:0] _T_389 = _T_385[3:2] | _T_385[1:0];
  wire [3:0] _T_393 = {_T_380,_T_384,_T_388,_T_389[1]};
  reg [5:0] nextAddr;
  wire [5:0] _T_400 = nextAddr + 6'h1;
  wire  _T_522 = ~_T_129;
  wire [5:0] _T_524 = _T_129 ? {{1'd0}, _T_150} : nextAddr;
  wire  _GEN_266 = 5'h0 == _T_524[4:0];
  wire  _GEN_0 = _GEN_266 | addresses_0_valid;
  wire  _GEN_267 = 5'h1 == _T_524[4:0];
  wire  _GEN_1 = _GEN_267 | addresses_1_valid;
  wire  _GEN_268 = 5'h2 == _T_524[4:0];
  wire  _GEN_2 = _GEN_268 | addresses_2_valid;
  wire  _GEN_269 = 5'h3 == _T_524[4:0];
  wire  _GEN_3 = _GEN_269 | addresses_3_valid;
  wire  _GEN_270 = 5'h4 == _T_524[4:0];
  wire  _GEN_4 = _GEN_270 | addresses_4_valid;
  wire  _GEN_271 = 5'h5 == _T_524[4:0];
  wire  _GEN_5 = _GEN_271 | addresses_5_valid;
  wire  _GEN_272 = 5'h6 == _T_524[4:0];
  wire  _GEN_6 = _GEN_272 | addresses_6_valid;
  wire  _GEN_273 = 5'h7 == _T_524[4:0];
  wire  _GEN_7 = _GEN_273 | addresses_7_valid;
  wire  _GEN_274 = 5'h8 == _T_524[4:0];
  wire  _GEN_8 = _GEN_274 | addresses_8_valid;
  wire  _GEN_275 = 5'h9 == _T_524[4:0];
  wire  _GEN_9 = _GEN_275 | addresses_9_valid;
  wire  _GEN_276 = 5'ha == _T_524[4:0];
  wire  _GEN_10 = _GEN_276 | addresses_10_valid;
  wire  _GEN_277 = 5'hb == _T_524[4:0];
  wire  _GEN_11 = _GEN_277 | addresses_11_valid;
  wire  _GEN_278 = 5'hc == _T_524[4:0];
  wire  _GEN_12 = _GEN_278 | addresses_12_valid;
  wire  _GEN_279 = 5'hd == _T_524[4:0];
  wire  _GEN_13 = _GEN_279 | addresses_13_valid;
  wire  _GEN_280 = 5'he == _T_524[4:0];
  wire  _GEN_14 = _GEN_280 | addresses_14_valid;
  wire  _GEN_281 = 5'hf == _T_524[4:0];
  wire  _GEN_15 = _GEN_281 | addresses_15_valid;
  wire  _GEN_282 = 5'h10 == _T_524[4:0];
  wire  _GEN_16 = _GEN_282 | addresses_16_valid;
  wire  _GEN_283 = 5'h11 == _T_524[4:0];
  wire  _GEN_17 = _GEN_283 | addresses_17_valid;
  wire  _GEN_284 = 5'h12 == _T_524[4:0];
  wire  _GEN_18 = _GEN_284 | addresses_18_valid;
  wire  _GEN_285 = 5'h13 == _T_524[4:0];
  wire  _GEN_19 = _GEN_285 | addresses_19_valid;
  wire  _GEN_286 = 5'h14 == _T_524[4:0];
  wire  _GEN_20 = _GEN_286 | addresses_20_valid;
  wire  _GEN_287 = 5'h15 == _T_524[4:0];
  wire  _GEN_21 = _GEN_287 | addresses_21_valid;
  wire  _GEN_288 = 5'h16 == _T_524[4:0];
  wire  _GEN_22 = _GEN_288 | addresses_22_valid;
  wire  _GEN_289 = 5'h17 == _T_524[4:0];
  wire  _GEN_23 = _GEN_289 | addresses_23_valid;
  wire  _GEN_290 = 5'h18 == _T_524[4:0];
  wire  _GEN_24 = _GEN_290 | addresses_24_valid;
  wire  _GEN_291 = 5'h19 == _T_524[4:0];
  wire  _GEN_25 = _GEN_291 | addresses_25_valid;
  wire  _GEN_292 = 5'h1a == _T_524[4:0];
  wire  _GEN_26 = _GEN_292 | addresses_26_valid;
  wire  _GEN_293 = 5'h1b == _T_524[4:0];
  wire  _GEN_27 = _GEN_293 | addresses_27_valid;
  wire  _GEN_294 = 5'h1c == _T_524[4:0];
  wire  _GEN_28 = _GEN_294 | addresses_28_valid;
  wire  _GEN_295 = 5'h1d == _T_524[4:0];
  wire  _GEN_29 = _GEN_295 | addresses_29_valid;
  wire  _GEN_296 = 5'h1e == _T_524[4:0];
  wire  _GEN_30 = _GEN_296 | addresses_30_valid;
  wire  _GEN_297 = 5'h1f == _T_524[4:0];
  wire  _GEN_31 = _GEN_297 | addresses_31_valid;
  wire [5:0] _T_531 = _T_522 ? _T_400 : nextAddr;
  wire  _T_532 = addresses_0_bits == io_w_1_addr;
  wire  _T_533 = addresses_0_valid & _T_532;
  wire  _T_534 = addresses_1_bits == io_w_1_addr;
  wire  _T_535 = addresses_1_valid & _T_534;
  wire  _T_536 = addresses_2_bits == io_w_1_addr;
  wire  _T_537 = addresses_2_valid & _T_536;
  wire  _T_538 = addresses_3_bits == io_w_1_addr;
  wire  _T_539 = addresses_3_valid & _T_538;
  wire  _T_540 = addresses_4_bits == io_w_1_addr;
  wire  _T_541 = addresses_4_valid & _T_540;
  wire  _T_542 = addresses_5_bits == io_w_1_addr;
  wire  _T_543 = addresses_5_valid & _T_542;
  wire  _T_544 = addresses_6_bits == io_w_1_addr;
  wire  _T_545 = addresses_6_valid & _T_544;
  wire  _T_546 = addresses_7_bits == io_w_1_addr;
  wire  _T_547 = addresses_7_valid & _T_546;
  wire  _T_548 = addresses_8_bits == io_w_1_addr;
  wire  _T_549 = addresses_8_valid & _T_548;
  wire  _T_550 = addresses_9_bits == io_w_1_addr;
  wire  _T_551 = addresses_9_valid & _T_550;
  wire  _T_552 = addresses_10_bits == io_w_1_addr;
  wire  _T_553 = addresses_10_valid & _T_552;
  wire  _T_554 = addresses_11_bits == io_w_1_addr;
  wire  _T_555 = addresses_11_valid & _T_554;
  wire  _T_556 = addresses_12_bits == io_w_1_addr;
  wire  _T_557 = addresses_12_valid & _T_556;
  wire  _T_558 = addresses_13_bits == io_w_1_addr;
  wire  _T_559 = addresses_13_valid & _T_558;
  wire  _T_560 = addresses_14_bits == io_w_1_addr;
  wire  _T_561 = addresses_14_valid & _T_560;
  wire  _T_562 = addresses_15_bits == io_w_1_addr;
  wire  _T_563 = addresses_15_valid & _T_562;
  wire  _T_564 = addresses_16_bits == io_w_1_addr;
  wire  _T_565 = addresses_16_valid & _T_564;
  wire  _T_566 = addresses_17_bits == io_w_1_addr;
  wire  _T_567 = addresses_17_valid & _T_566;
  wire  _T_568 = addresses_18_bits == io_w_1_addr;
  wire  _T_569 = addresses_18_valid & _T_568;
  wire  _T_570 = addresses_19_bits == io_w_1_addr;
  wire  _T_571 = addresses_19_valid & _T_570;
  wire  _T_572 = addresses_20_bits == io_w_1_addr;
  wire  _T_573 = addresses_20_valid & _T_572;
  wire  _T_574 = addresses_21_bits == io_w_1_addr;
  wire  _T_575 = addresses_21_valid & _T_574;
  wire  _T_576 = addresses_22_bits == io_w_1_addr;
  wire  _T_577 = addresses_22_valid & _T_576;
  wire  _T_578 = addresses_23_bits == io_w_1_addr;
  wire  _T_579 = addresses_23_valid & _T_578;
  wire  _T_580 = addresses_24_bits == io_w_1_addr;
  wire  _T_581 = addresses_24_valid & _T_580;
  wire  _T_582 = addresses_25_bits == io_w_1_addr;
  wire  _T_583 = addresses_25_valid & _T_582;
  wire  _T_584 = addresses_26_bits == io_w_1_addr;
  wire  _T_585 = addresses_26_valid & _T_584;
  wire  _T_586 = addresses_27_bits == io_w_1_addr;
  wire  _T_587 = addresses_27_valid & _T_586;
  wire  _T_588 = addresses_28_bits == io_w_1_addr;
  wire  _T_589 = addresses_28_valid & _T_588;
  wire  _T_590 = addresses_29_bits == io_w_1_addr;
  wire  _T_591 = addresses_29_valid & _T_590;
  wire  _T_592 = addresses_30_bits == io_w_1_addr;
  wire  _T_593 = addresses_30_valid & _T_592;
  wire  _T_594 = addresses_31_bits == io_w_1_addr;
  wire  _T_595 = addresses_31_valid & _T_594;
  wire [7:0] _T_603 = {_T_547,_T_545,_T_543,_T_541,_T_539,_T_537,_T_535,_T_533};
  wire [15:0] _T_611 = {_T_563,_T_561,_T_559,_T_557,_T_555,_T_553,_T_551,_T_549,_T_603};
  wire [7:0] _T_618 = {_T_579,_T_577,_T_575,_T_573,_T_571,_T_569,_T_567,_T_565};
  wire [31:0] _T_627 = {_T_595,_T_593,_T_591,_T_589,_T_587,_T_585,_T_583,_T_581,_T_618,_T_611};
  wire  _T_628 = _T_627 != 32'h0;
  wire  _T_631 = |_T_627[31:16];
  wire [15:0] _T_632 = _T_627[31:16] | _T_627[15:0];
  wire  _T_635 = |_T_632[15:8];
  wire [7:0] _T_636 = _T_632[15:8] | _T_632[7:0];
  wire  _T_639 = |_T_636[7:4];
  wire [3:0] _T_640 = _T_636[7:4] | _T_636[3:0];
  wire  _T_643 = |_T_640[3:2];
  wire [1:0] _T_644 = _T_640[3:2] | _T_640[1:0];
  wire [4:0] _T_649 = {_T_631,_T_635,_T_639,_T_643,_T_644[1]};
  wire  _T_650 = ~_T_628;
  wire  _T_651 = io_w_1_en & _T_650;
  wire [5:0] _T_652 = _T_628 ? {{1'd0}, _T_649} : _T_531;
  wire  _GEN_298 = 5'h0 == _T_652[4:0];
  wire  _GEN_133 = _GEN_298 | _GEN_0;
  wire  _GEN_299 = 5'h1 == _T_652[4:0];
  wire  _GEN_134 = _GEN_299 | _GEN_1;
  wire  _GEN_300 = 5'h2 == _T_652[4:0];
  wire  _GEN_135 = _GEN_300 | _GEN_2;
  wire  _GEN_301 = 5'h3 == _T_652[4:0];
  wire  _GEN_136 = _GEN_301 | _GEN_3;
  wire  _GEN_302 = 5'h4 == _T_652[4:0];
  wire  _GEN_137 = _GEN_302 | _GEN_4;
  wire  _GEN_303 = 5'h5 == _T_652[4:0];
  wire  _GEN_138 = _GEN_303 | _GEN_5;
  wire  _GEN_304 = 5'h6 == _T_652[4:0];
  wire  _GEN_139 = _GEN_304 | _GEN_6;
  wire  _GEN_305 = 5'h7 == _T_652[4:0];
  wire  _GEN_140 = _GEN_305 | _GEN_7;
  wire  _GEN_306 = 5'h8 == _T_652[4:0];
  wire  _GEN_141 = _GEN_306 | _GEN_8;
  wire  _GEN_307 = 5'h9 == _T_652[4:0];
  wire  _GEN_142 = _GEN_307 | _GEN_9;
  wire  _GEN_308 = 5'ha == _T_652[4:0];
  wire  _GEN_143 = _GEN_308 | _GEN_10;
  wire  _GEN_309 = 5'hb == _T_652[4:0];
  wire  _GEN_144 = _GEN_309 | _GEN_11;
  wire  _GEN_310 = 5'hc == _T_652[4:0];
  wire  _GEN_145 = _GEN_310 | _GEN_12;
  wire  _GEN_311 = 5'hd == _T_652[4:0];
  wire  _GEN_146 = _GEN_311 | _GEN_13;
  wire  _GEN_312 = 5'he == _T_652[4:0];
  wire  _GEN_147 = _GEN_312 | _GEN_14;
  wire  _GEN_313 = 5'hf == _T_652[4:0];
  wire  _GEN_148 = _GEN_313 | _GEN_15;
  wire  _GEN_314 = 5'h10 == _T_652[4:0];
  wire  _GEN_149 = _GEN_314 | _GEN_16;
  wire  _GEN_315 = 5'h11 == _T_652[4:0];
  wire  _GEN_150 = _GEN_315 | _GEN_17;
  wire  _GEN_316 = 5'h12 == _T_652[4:0];
  wire  _GEN_151 = _GEN_316 | _GEN_18;
  wire  _GEN_317 = 5'h13 == _T_652[4:0];
  wire  _GEN_152 = _GEN_317 | _GEN_19;
  wire  _GEN_318 = 5'h14 == _T_652[4:0];
  wire  _GEN_153 = _GEN_318 | _GEN_20;
  wire  _GEN_319 = 5'h15 == _T_652[4:0];
  wire  _GEN_154 = _GEN_319 | _GEN_21;
  wire  _GEN_320 = 5'h16 == _T_652[4:0];
  wire  _GEN_155 = _GEN_320 | _GEN_22;
  wire  _GEN_321 = 5'h17 == _T_652[4:0];
  wire  _GEN_156 = _GEN_321 | _GEN_23;
  wire  _GEN_322 = 5'h18 == _T_652[4:0];
  wire  _GEN_157 = _GEN_322 | _GEN_24;
  wire  _GEN_323 = 5'h19 == _T_652[4:0];
  wire  _GEN_158 = _GEN_323 | _GEN_25;
  wire  _GEN_324 = 5'h1a == _T_652[4:0];
  wire  _GEN_159 = _GEN_324 | _GEN_26;
  wire  _GEN_325 = 5'h1b == _T_652[4:0];
  wire  _GEN_160 = _GEN_325 | _GEN_27;
  wire  _GEN_326 = 5'h1c == _T_652[4:0];
  wire  _GEN_161 = _GEN_326 | _GEN_28;
  wire  _GEN_327 = 5'h1d == _T_652[4:0];
  wire  _GEN_162 = _GEN_327 | _GEN_29;
  wire  _GEN_328 = 5'h1e == _T_652[4:0];
  wire  _GEN_163 = _GEN_328 | _GEN_30;
  wire  _GEN_329 = 5'h1f == _T_652[4:0];
  wire  _GEN_164 = _GEN_329 | _GEN_31;
  wire [5:0] _T_658 = _T_531 + 6'h1;
  wire [5:0] nextAddrUpdate = _T_651 ? _T_658 : _T_531;
  wire  _T_659 = nextAddrUpdate <= 6'h20;
  wire  _T_661 = _T_659 | reset;
  wire  _T_662 = ~_T_661;
  assign mem__T_152_addr = {_T_132,_T_149};
  assign mem__T_152_data = mem[mem__T_152_addr];
  assign mem__T_274_addr = {_T_254,_T_271};
  assign mem__T_274_data = mem[mem__T_274_addr];
  assign mem__T_396_addr = {_T_376,_T_393};
  assign mem__T_396_data = mem[mem__T_396_addr];
  assign mem__T_528_data = 32'h0;
  assign mem__T_528_addr = _T_524[4:0];
  assign mem__T_528_mask = 1'h1;
  assign mem__T_528_en = 1'h1;
  assign mem__T_656_data = io_w_1_data;
  assign mem__T_656_addr = _T_652[4:0];
  assign mem__T_656_mask = 1'h1;
  assign mem__T_656_en = io_w_1_en;
  assign io_r_1_data = _T_251 ? mem__T_274_data : 32'h0;
  assign io_r_2_data = _T_373 ? mem__T_396_data : 32'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  addresses_0_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  addresses_0_bits = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  addresses_1_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  addresses_1_bits = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  addresses_2_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  addresses_2_bits = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  addresses_3_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  addresses_3_bits = _RAND_8[4:0];
  _RAND_9 = {1{`RANDOM}};
  addresses_4_valid = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  addresses_4_bits = _RAND_10[4:0];
  _RAND_11 = {1{`RANDOM}};
  addresses_5_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  addresses_5_bits = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  addresses_6_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  addresses_6_bits = _RAND_14[4:0];
  _RAND_15 = {1{`RANDOM}};
  addresses_7_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  addresses_7_bits = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  addresses_8_valid = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  addresses_8_bits = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  addresses_9_valid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  addresses_9_bits = _RAND_20[4:0];
  _RAND_21 = {1{`RANDOM}};
  addresses_10_valid = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  addresses_10_bits = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  addresses_11_valid = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  addresses_11_bits = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  addresses_12_valid = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  addresses_12_bits = _RAND_26[4:0];
  _RAND_27 = {1{`RANDOM}};
  addresses_13_valid = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  addresses_13_bits = _RAND_28[4:0];
  _RAND_29 = {1{`RANDOM}};
  addresses_14_valid = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  addresses_14_bits = _RAND_30[4:0];
  _RAND_31 = {1{`RANDOM}};
  addresses_15_valid = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  addresses_15_bits = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  addresses_16_valid = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  addresses_16_bits = _RAND_34[4:0];
  _RAND_35 = {1{`RANDOM}};
  addresses_17_valid = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  addresses_17_bits = _RAND_36[4:0];
  _RAND_37 = {1{`RANDOM}};
  addresses_18_valid = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  addresses_18_bits = _RAND_38[4:0];
  _RAND_39 = {1{`RANDOM}};
  addresses_19_valid = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  addresses_19_bits = _RAND_40[4:0];
  _RAND_41 = {1{`RANDOM}};
  addresses_20_valid = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  addresses_20_bits = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  addresses_21_valid = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  addresses_21_bits = _RAND_44[4:0];
  _RAND_45 = {1{`RANDOM}};
  addresses_22_valid = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  addresses_22_bits = _RAND_46[4:0];
  _RAND_47 = {1{`RANDOM}};
  addresses_23_valid = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  addresses_23_bits = _RAND_48[4:0];
  _RAND_49 = {1{`RANDOM}};
  addresses_24_valid = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  addresses_24_bits = _RAND_50[4:0];
  _RAND_51 = {1{`RANDOM}};
  addresses_25_valid = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  addresses_25_bits = _RAND_52[4:0];
  _RAND_53 = {1{`RANDOM}};
  addresses_26_valid = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  addresses_26_bits = _RAND_54[4:0];
  _RAND_55 = {1{`RANDOM}};
  addresses_27_valid = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  addresses_27_bits = _RAND_56[4:0];
  _RAND_57 = {1{`RANDOM}};
  addresses_28_valid = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  addresses_28_bits = _RAND_58[4:0];
  _RAND_59 = {1{`RANDOM}};
  addresses_29_valid = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  addresses_29_bits = _RAND_60[4:0];
  _RAND_61 = {1{`RANDOM}};
  addresses_30_valid = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  addresses_30_bits = _RAND_62[4:0];
  _RAND_63 = {1{`RANDOM}};
  addresses_31_valid = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  addresses_31_bits = _RAND_64[4:0];
  _RAND_65 = {1{`RANDOM}};
  nextAddr = _RAND_65[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_528_en & mem__T_528_mask) begin
      mem[mem__T_528_addr] <= mem__T_528_data;
    end
    if(mem__T_656_en & mem__T_656_mask) begin
      mem[mem__T_656_addr] <= mem__T_656_data;
    end
    if (metaReset) begin
      addresses_0_valid <= 1'h0;
    end else if (reset) begin
      addresses_0_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_0_valid <= _GEN_133;
    end else begin
      addresses_0_valid <= _GEN_0;
    end
    if (metaReset) begin
      addresses_0_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h0 == _T_652[4:0]) begin
        addresses_0_bits <= io_w_1_addr;
      end else if (5'h0 == _T_524[4:0]) begin
        addresses_0_bits <= 5'h0;
      end
    end else if (5'h0 == _T_524[4:0]) begin
      addresses_0_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_1_valid <= 1'h0;
    end else if (reset) begin
      addresses_1_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_1_valid <= _GEN_134;
    end else begin
      addresses_1_valid <= _GEN_1;
    end
    if (metaReset) begin
      addresses_1_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h1 == _T_652[4:0]) begin
        addresses_1_bits <= io_w_1_addr;
      end else if (5'h1 == _T_524[4:0]) begin
        addresses_1_bits <= 5'h0;
      end
    end else if (5'h1 == _T_524[4:0]) begin
      addresses_1_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_2_valid <= 1'h0;
    end else if (reset) begin
      addresses_2_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_2_valid <= _GEN_135;
    end else begin
      addresses_2_valid <= _GEN_2;
    end
    if (metaReset) begin
      addresses_2_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h2 == _T_652[4:0]) begin
        addresses_2_bits <= io_w_1_addr;
      end else if (5'h2 == _T_524[4:0]) begin
        addresses_2_bits <= 5'h0;
      end
    end else if (5'h2 == _T_524[4:0]) begin
      addresses_2_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_3_valid <= 1'h0;
    end else if (reset) begin
      addresses_3_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_3_valid <= _GEN_136;
    end else begin
      addresses_3_valid <= _GEN_3;
    end
    if (metaReset) begin
      addresses_3_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h3 == _T_652[4:0]) begin
        addresses_3_bits <= io_w_1_addr;
      end else if (5'h3 == _T_524[4:0]) begin
        addresses_3_bits <= 5'h0;
      end
    end else if (5'h3 == _T_524[4:0]) begin
      addresses_3_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_4_valid <= 1'h0;
    end else if (reset) begin
      addresses_4_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_4_valid <= _GEN_137;
    end else begin
      addresses_4_valid <= _GEN_4;
    end
    if (metaReset) begin
      addresses_4_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h4 == _T_652[4:0]) begin
        addresses_4_bits <= io_w_1_addr;
      end else if (5'h4 == _T_524[4:0]) begin
        addresses_4_bits <= 5'h0;
      end
    end else if (5'h4 == _T_524[4:0]) begin
      addresses_4_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_5_valid <= 1'h0;
    end else if (reset) begin
      addresses_5_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_5_valid <= _GEN_138;
    end else begin
      addresses_5_valid <= _GEN_5;
    end
    if (metaReset) begin
      addresses_5_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h5 == _T_652[4:0]) begin
        addresses_5_bits <= io_w_1_addr;
      end else if (5'h5 == _T_524[4:0]) begin
        addresses_5_bits <= 5'h0;
      end
    end else if (5'h5 == _T_524[4:0]) begin
      addresses_5_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_6_valid <= 1'h0;
    end else if (reset) begin
      addresses_6_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_6_valid <= _GEN_139;
    end else begin
      addresses_6_valid <= _GEN_6;
    end
    if (metaReset) begin
      addresses_6_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h6 == _T_652[4:0]) begin
        addresses_6_bits <= io_w_1_addr;
      end else if (5'h6 == _T_524[4:0]) begin
        addresses_6_bits <= 5'h0;
      end
    end else if (5'h6 == _T_524[4:0]) begin
      addresses_6_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_7_valid <= 1'h0;
    end else if (reset) begin
      addresses_7_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_7_valid <= _GEN_140;
    end else begin
      addresses_7_valid <= _GEN_7;
    end
    if (metaReset) begin
      addresses_7_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h7 == _T_652[4:0]) begin
        addresses_7_bits <= io_w_1_addr;
      end else if (5'h7 == _T_524[4:0]) begin
        addresses_7_bits <= 5'h0;
      end
    end else if (5'h7 == _T_524[4:0]) begin
      addresses_7_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_8_valid <= 1'h0;
    end else if (reset) begin
      addresses_8_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_8_valid <= _GEN_141;
    end else begin
      addresses_8_valid <= _GEN_8;
    end
    if (metaReset) begin
      addresses_8_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h8 == _T_652[4:0]) begin
        addresses_8_bits <= io_w_1_addr;
      end else if (5'h8 == _T_524[4:0]) begin
        addresses_8_bits <= 5'h0;
      end
    end else if (5'h8 == _T_524[4:0]) begin
      addresses_8_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_9_valid <= 1'h0;
    end else if (reset) begin
      addresses_9_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_9_valid <= _GEN_142;
    end else begin
      addresses_9_valid <= _GEN_9;
    end
    if (metaReset) begin
      addresses_9_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h9 == _T_652[4:0]) begin
        addresses_9_bits <= io_w_1_addr;
      end else if (5'h9 == _T_524[4:0]) begin
        addresses_9_bits <= 5'h0;
      end
    end else if (5'h9 == _T_524[4:0]) begin
      addresses_9_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_10_valid <= 1'h0;
    end else if (reset) begin
      addresses_10_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_10_valid <= _GEN_143;
    end else begin
      addresses_10_valid <= _GEN_10;
    end
    if (metaReset) begin
      addresses_10_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'ha == _T_652[4:0]) begin
        addresses_10_bits <= io_w_1_addr;
      end else if (5'ha == _T_524[4:0]) begin
        addresses_10_bits <= 5'h0;
      end
    end else if (5'ha == _T_524[4:0]) begin
      addresses_10_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_11_valid <= 1'h0;
    end else if (reset) begin
      addresses_11_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_11_valid <= _GEN_144;
    end else begin
      addresses_11_valid <= _GEN_11;
    end
    if (metaReset) begin
      addresses_11_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'hb == _T_652[4:0]) begin
        addresses_11_bits <= io_w_1_addr;
      end else if (5'hb == _T_524[4:0]) begin
        addresses_11_bits <= 5'h0;
      end
    end else if (5'hb == _T_524[4:0]) begin
      addresses_11_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_12_valid <= 1'h0;
    end else if (reset) begin
      addresses_12_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_12_valid <= _GEN_145;
    end else begin
      addresses_12_valid <= _GEN_12;
    end
    if (metaReset) begin
      addresses_12_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'hc == _T_652[4:0]) begin
        addresses_12_bits <= io_w_1_addr;
      end else if (5'hc == _T_524[4:0]) begin
        addresses_12_bits <= 5'h0;
      end
    end else if (5'hc == _T_524[4:0]) begin
      addresses_12_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_13_valid <= 1'h0;
    end else if (reset) begin
      addresses_13_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_13_valid <= _GEN_146;
    end else begin
      addresses_13_valid <= _GEN_13;
    end
    if (metaReset) begin
      addresses_13_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'hd == _T_652[4:0]) begin
        addresses_13_bits <= io_w_1_addr;
      end else if (5'hd == _T_524[4:0]) begin
        addresses_13_bits <= 5'h0;
      end
    end else if (5'hd == _T_524[4:0]) begin
      addresses_13_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_14_valid <= 1'h0;
    end else if (reset) begin
      addresses_14_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_14_valid <= _GEN_147;
    end else begin
      addresses_14_valid <= _GEN_14;
    end
    if (metaReset) begin
      addresses_14_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'he == _T_652[4:0]) begin
        addresses_14_bits <= io_w_1_addr;
      end else if (5'he == _T_524[4:0]) begin
        addresses_14_bits <= 5'h0;
      end
    end else if (5'he == _T_524[4:0]) begin
      addresses_14_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_15_valid <= 1'h0;
    end else if (reset) begin
      addresses_15_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_15_valid <= _GEN_148;
    end else begin
      addresses_15_valid <= _GEN_15;
    end
    if (metaReset) begin
      addresses_15_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'hf == _T_652[4:0]) begin
        addresses_15_bits <= io_w_1_addr;
      end else if (5'hf == _T_524[4:0]) begin
        addresses_15_bits <= 5'h0;
      end
    end else if (5'hf == _T_524[4:0]) begin
      addresses_15_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_16_valid <= 1'h0;
    end else if (reset) begin
      addresses_16_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_16_valid <= _GEN_149;
    end else begin
      addresses_16_valid <= _GEN_16;
    end
    if (metaReset) begin
      addresses_16_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h10 == _T_652[4:0]) begin
        addresses_16_bits <= io_w_1_addr;
      end else if (5'h10 == _T_524[4:0]) begin
        addresses_16_bits <= 5'h0;
      end
    end else if (5'h10 == _T_524[4:0]) begin
      addresses_16_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_17_valid <= 1'h0;
    end else if (reset) begin
      addresses_17_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_17_valid <= _GEN_150;
    end else begin
      addresses_17_valid <= _GEN_17;
    end
    if (metaReset) begin
      addresses_17_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h11 == _T_652[4:0]) begin
        addresses_17_bits <= io_w_1_addr;
      end else if (5'h11 == _T_524[4:0]) begin
        addresses_17_bits <= 5'h0;
      end
    end else if (5'h11 == _T_524[4:0]) begin
      addresses_17_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_18_valid <= 1'h0;
    end else if (reset) begin
      addresses_18_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_18_valid <= _GEN_151;
    end else begin
      addresses_18_valid <= _GEN_18;
    end
    if (metaReset) begin
      addresses_18_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h12 == _T_652[4:0]) begin
        addresses_18_bits <= io_w_1_addr;
      end else if (5'h12 == _T_524[4:0]) begin
        addresses_18_bits <= 5'h0;
      end
    end else if (5'h12 == _T_524[4:0]) begin
      addresses_18_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_19_valid <= 1'h0;
    end else if (reset) begin
      addresses_19_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_19_valid <= _GEN_152;
    end else begin
      addresses_19_valid <= _GEN_19;
    end
    if (metaReset) begin
      addresses_19_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h13 == _T_652[4:0]) begin
        addresses_19_bits <= io_w_1_addr;
      end else if (5'h13 == _T_524[4:0]) begin
        addresses_19_bits <= 5'h0;
      end
    end else if (5'h13 == _T_524[4:0]) begin
      addresses_19_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_20_valid <= 1'h0;
    end else if (reset) begin
      addresses_20_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_20_valid <= _GEN_153;
    end else begin
      addresses_20_valid <= _GEN_20;
    end
    if (metaReset) begin
      addresses_20_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h14 == _T_652[4:0]) begin
        addresses_20_bits <= io_w_1_addr;
      end else if (5'h14 == _T_524[4:0]) begin
        addresses_20_bits <= 5'h0;
      end
    end else if (5'h14 == _T_524[4:0]) begin
      addresses_20_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_21_valid <= 1'h0;
    end else if (reset) begin
      addresses_21_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_21_valid <= _GEN_154;
    end else begin
      addresses_21_valid <= _GEN_21;
    end
    if (metaReset) begin
      addresses_21_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h15 == _T_652[4:0]) begin
        addresses_21_bits <= io_w_1_addr;
      end else if (5'h15 == _T_524[4:0]) begin
        addresses_21_bits <= 5'h0;
      end
    end else if (5'h15 == _T_524[4:0]) begin
      addresses_21_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_22_valid <= 1'h0;
    end else if (reset) begin
      addresses_22_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_22_valid <= _GEN_155;
    end else begin
      addresses_22_valid <= _GEN_22;
    end
    if (metaReset) begin
      addresses_22_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h16 == _T_652[4:0]) begin
        addresses_22_bits <= io_w_1_addr;
      end else if (5'h16 == _T_524[4:0]) begin
        addresses_22_bits <= 5'h0;
      end
    end else if (5'h16 == _T_524[4:0]) begin
      addresses_22_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_23_valid <= 1'h0;
    end else if (reset) begin
      addresses_23_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_23_valid <= _GEN_156;
    end else begin
      addresses_23_valid <= _GEN_23;
    end
    if (metaReset) begin
      addresses_23_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h17 == _T_652[4:0]) begin
        addresses_23_bits <= io_w_1_addr;
      end else if (5'h17 == _T_524[4:0]) begin
        addresses_23_bits <= 5'h0;
      end
    end else if (5'h17 == _T_524[4:0]) begin
      addresses_23_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_24_valid <= 1'h0;
    end else if (reset) begin
      addresses_24_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_24_valid <= _GEN_157;
    end else begin
      addresses_24_valid <= _GEN_24;
    end
    if (metaReset) begin
      addresses_24_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h18 == _T_652[4:0]) begin
        addresses_24_bits <= io_w_1_addr;
      end else if (5'h18 == _T_524[4:0]) begin
        addresses_24_bits <= 5'h0;
      end
    end else if (5'h18 == _T_524[4:0]) begin
      addresses_24_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_25_valid <= 1'h0;
    end else if (reset) begin
      addresses_25_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_25_valid <= _GEN_158;
    end else begin
      addresses_25_valid <= _GEN_25;
    end
    if (metaReset) begin
      addresses_25_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h19 == _T_652[4:0]) begin
        addresses_25_bits <= io_w_1_addr;
      end else if (5'h19 == _T_524[4:0]) begin
        addresses_25_bits <= 5'h0;
      end
    end else if (5'h19 == _T_524[4:0]) begin
      addresses_25_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_26_valid <= 1'h0;
    end else if (reset) begin
      addresses_26_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_26_valid <= _GEN_159;
    end else begin
      addresses_26_valid <= _GEN_26;
    end
    if (metaReset) begin
      addresses_26_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h1a == _T_652[4:0]) begin
        addresses_26_bits <= io_w_1_addr;
      end else if (5'h1a == _T_524[4:0]) begin
        addresses_26_bits <= 5'h0;
      end
    end else if (5'h1a == _T_524[4:0]) begin
      addresses_26_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_27_valid <= 1'h0;
    end else if (reset) begin
      addresses_27_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_27_valid <= _GEN_160;
    end else begin
      addresses_27_valid <= _GEN_27;
    end
    if (metaReset) begin
      addresses_27_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h1b == _T_652[4:0]) begin
        addresses_27_bits <= io_w_1_addr;
      end else if (5'h1b == _T_524[4:0]) begin
        addresses_27_bits <= 5'h0;
      end
    end else if (5'h1b == _T_524[4:0]) begin
      addresses_27_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_28_valid <= 1'h0;
    end else if (reset) begin
      addresses_28_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_28_valid <= _GEN_161;
    end else begin
      addresses_28_valid <= _GEN_28;
    end
    if (metaReset) begin
      addresses_28_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h1c == _T_652[4:0]) begin
        addresses_28_bits <= io_w_1_addr;
      end else if (5'h1c == _T_524[4:0]) begin
        addresses_28_bits <= 5'h0;
      end
    end else if (5'h1c == _T_524[4:0]) begin
      addresses_28_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_29_valid <= 1'h0;
    end else if (reset) begin
      addresses_29_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_29_valid <= _GEN_162;
    end else begin
      addresses_29_valid <= _GEN_29;
    end
    if (metaReset) begin
      addresses_29_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h1d == _T_652[4:0]) begin
        addresses_29_bits <= io_w_1_addr;
      end else if (5'h1d == _T_524[4:0]) begin
        addresses_29_bits <= 5'h0;
      end
    end else if (5'h1d == _T_524[4:0]) begin
      addresses_29_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_30_valid <= 1'h0;
    end else if (reset) begin
      addresses_30_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_30_valid <= _GEN_163;
    end else begin
      addresses_30_valid <= _GEN_30;
    end
    if (metaReset) begin
      addresses_30_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h1e == _T_652[4:0]) begin
        addresses_30_bits <= io_w_1_addr;
      end else if (5'h1e == _T_524[4:0]) begin
        addresses_30_bits <= 5'h0;
      end
    end else if (5'h1e == _T_524[4:0]) begin
      addresses_30_bits <= 5'h0;
    end
    if (metaReset) begin
      addresses_31_valid <= 1'h0;
    end else if (reset) begin
      addresses_31_valid <= 1'h0;
    end else if (io_w_1_en) begin
      addresses_31_valid <= _GEN_164;
    end else begin
      addresses_31_valid <= _GEN_31;
    end
    if (metaReset) begin
      addresses_31_bits <= 5'h0;
    end else if (io_w_1_en) begin
      if (5'h1f == _T_652[4:0]) begin
        addresses_31_bits <= io_w_1_addr;
      end else if (5'h1f == _T_524[4:0]) begin
        addresses_31_bits <= 5'h0;
      end
    end else if (5'h1f == _T_524[4:0]) begin
      addresses_31_bits <= 5'h0;
    end
    if (metaReset) begin
      nextAddr <= 6'h0;
    end else if (reset) begin
      nextAddr <= 6'h0;
    end else if (_T_651) begin
      nextAddr <= _T_658;
    end else if (_T_522) begin
      nextAddr <= _T_400;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_662) begin
          $fwrite(32'h80000002,"Assertion failed: SparseMem ran out of space with size %d, increase size in ReplaceMemsTransform!\n    at SparseMem.scala:102 assert(nextAddrUpdate <= depth.U,\n",6'h20);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_662) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Core(
  input         metaReset,
  input         clock,
  input         reset,
  output [31:0] io_imem_req_bits_addr,
  input  [31:0] io_imem_resp_bits_data,
  output [31:0] io_dmem_req_bits_addr,
  output [31:0] io_dmem_req_bits_data,
  output        io_dmem_req_bits_fcn,
  output [2:0]  io_dmem_req_bits_typ,
  input  [31:0] io_dmem_resp_bits_data,
  output        _GEN_411,
  output        _GEN_405,
  output        _GEN_92,
  output        _GEN_52,
  output        _GEN_305,
  output        _GEN_200,
  output        _GEN_149,
  output        _GEN_426,
  output        _GEN_291,
  output        _GEN_1_0,
  output        _GEN_25,
  output        _GEN_248,
  output        _GEN_107,
  output        _GEN_134,
  output        _GEN_206,
  output        _GEN_40,
  output        _GEN_306,
  output        _GEN_233,
  output        _GEN_128,
  output        _GEN_384,
  output        _GEN_191,
  output        _GEN_16,
  output        _GEN_227,
  output        _GEN_19,
  output        _GEN_327,
  output        _GEN_113,
  output        _GEN_46,
  output        _GEN_299,
  output        _GEN_390,
  output        _GEN_73,
  output        _GEN_212,
  output        _GEN_10,
  output        _GEN_285,
  output        _GEN_318,
  output        _GEN_312,
  output        _GEN_31,
  output        _GEN_311,
  output        _GEN_67,
  output        _GEN_320,
  output        _GEN_399,
  output        _GEN_215,
  output        _GEN_221,
  output        _GEN_101,
  output        _GEN_110,
  output        _GEN_387,
  output        _GEN_283,
  output        _GEN_314,
  output        _GEN_178,
  output        _GEN_209,
  output        _GEN_300,
  output        _GEN_279,
  output        _GEN_269,
  output        _GEN_28,
  output        _GEN_277,
  output        _GEN_378,
  output        _GEN_368,
  output        _GEN_55,
  output        _GEN_377,
  output        _GEN_194,
  output        _GEN_22,
  output        _GEN_12,
  output        _GEN_294,
  output        _GEN_13,
  output        _GEN_49,
  output        _GEN_116,
  output        _GEN_393,
  output        _GEN_362,
  output        _GEN_7,
  output        _GEN_461,
  output        _GEN_34,
  output        _GEN_122,
  output        _GEN_308,
  output        _GEN_263,
  output        _GEN_95,
  output        _GEN_230,
  output        _GEN_293,
  output        _GEN_184,
  output        _GEN_1_1,
  output        _GEN_10_0,
  output        _GEN_197,
  output        _GEN_187,
  output        _GEN_449,
  output        _GEN_288,
  output        _GEN_104,
  output        _GEN_265,
  output        _GEN_296,
  output        _GEN_160,
  output        _GEN_172,
  output        _GEN_203,
  output        _GEN_245,
  output        _GEN_0,
  output        _GEN_272,
  output        _GEN_271,
  output        _GEN_37,
  output        _GEN_166,
  output        _GEN_280,
  output        _GEN_286,
  output        _GEN_381,
  output        _GEN_371,
  output        _GEN_266,
  output        _GEN_16_0,
  output        _GEN_22_0,
  output        _GEN_302,
  output        _GEN_344,
  output        _GEN_282,
  output        _GEN_443,
  output        _GEN_16_1,
  output        _GEN_251,
  output        _GEN_10_1,
  output        _GEN_259,
  output        _GEN_98,
  output        _GEN_6,
  output        _GEN_350,
  output        _GEN_365,
  output        _GEN_15,
  output        _GEN_152,
  output        _GEN_446,
  output        _GEN_332,
  output        _GEN_326,
  output        _GEN_19_0,
  output        _GEN_148,
  output        _GEN_359,
  output        _GEN_15_0,
  output        _GEN_87,
  output        _GEN_458,
  output        _GEN_452,
  output        _GEN_13_0,
  output        _GEN_3,
  output        _GEN_347,
  output        _GEN_274,
  output        _GEN_425,
  output        _GEN_239,
  output        _GEN_232,
  output        _GEN_190,
  output        _GEN_154,
  output        _GEN_289,
  output        _GEN_431,
  output        _GEN_181,
  output        _GEN_253,
  output        _GEN_254,
  output        _GEN_353,
  output        _GEN_72,
  output        _GEN_175,
  output        _GEN_169,
  output        _GEN_260,
  output        _GEN_4_0,
  output        _GEN_275,
  output        _GEN_247,
  output        _GEN_268,
  output        _GEN_9,
  output        _GEN_338,
  output        _GEN_374,
  output        _GEN_242,
  output        _GEN_214,
  output        _GEN_250,
  output        _GEN_455,
  output        _GEN_241,
  output        _GEN_142,
  output        _GEN_136,
  output        _GEN_413,
  output        _GEN_235,
  output        _GEN_236,
  output        _GEN_262,
  output        _GEN_335,
  output        _GEN_54,
  output        _GEN_313,
  output        _GEN_18,
  output        _GEN_69,
  output        _GEN_157,
  output        _GEN_434,
  output        _GEN_248_0,
  output        _GEN_257,
  output        _GEN_320_0,
  output        _GEN_75,
  output        _GEN_356,
  output        _GEN_12_0,
  output        _GEN_90,
  output        _GEN_163,
  output        _GEN_419,
  output        _GEN_314_0,
  output        _GEN_7_0,
  output        _GEN_130,
  output        _GEN_341,
  output        _GEN_440,
  output        _GEN_229,
  output        _GEN_299_0,
  output        _GEN_121,
  output        _GEN_256,
  output        _GEN_398,
  output        _GEN_81,
  output        _GEN_407,
  output        _GEN_149_0,
  output        _GEN_416,
  output        _GEN_281,
  output        _GEN_15_1,
  output        _GEN_380,
  output        _GEN_57,
  output        _GEN_145,
  output        _GEN_296_0,
  output        _GEN_223,
  output        _GEN_118,
  output        _GEN_322,
  output        _GEN_422,
  output        _GEN_244,
  output        _GEN_124,
  output        _GEN_103,
  output        _GEN_238,
  output        _GEN_329,
  output        _GEN_63,
  output        _GEN_151,
  output        _GEN_202,
  output        _GEN_6_0,
  output        _GEN_196,
  output        _GEN_437,
  output        _GEN_302_0,
  output        _GEN_295,
  output        _GEN_301,
  output        _GEN_310,
  output        _GEN_401,
  output        _GEN_395,
  output        _GEN_78,
  output        _GEN_84,
  output        _GEN_217,
  output        _GEN_428,
  output        _GEN_308_0,
  output        _GEN_323,
  output        _GEN_36,
  output        _GEN_42,
  output        _GEN_317,
  output        _GEN_316,
  output        _GEN_139,
  output        _GEN_404,
  output        _GEN_290,
  output        _GEN_18_0,
  output        _GEN_226,
  output        _GEN_106,
  output        _GEN_51,
  output        _GEN_45,
  output        _GEN_9_0,
  output        _GEN_367,
  output        _GEN_319,
  output        _GEN_284,
  output        _GEN_274_0,
  output        _GEN_39,
  output        _GEN_383,
  output        _GEN_373,
  output        _GEN_66,
  output        _GEN_18_1,
  output        _GEN_410,
  output        _GEN_24,
  output        _GEN_305_0,
  output        _GEN_112,
  output        _GEN_211,
  output        _GEN_220,
  output        _GEN_8,
  output        _GEN_2,
  output        _GEN_311_0,
  output        _GEN_133,
  output        _GEN_127,
  output        _GEN_288_0,
  output        _GEN_389,
  output        _GEN_91,
  output        _GEN_205,
  output        _GEN_100,
  output        _GEN_304,
  output        _GEN_60,
  output        _GEN_298,
  output        _GEN_189,
  output        _GEN_199,
  output        _GEN_177,
  output        _GEN_12_1,
  output        _GEN_268_0,
  output        _GEN_94,
  output        _GEN_376,
  output        _GEN_162,
  output        _GEN_193,
  output        _GEN_208,
  output        _GEN_454,
  output        _GEN_293_0,
  output        _GEN_261,
  output        _GEN_115,
  output        _GEN_27,
  output        _GEN_270,
  output        _GEN_392,
  output        _GEN_361,
  output        _GEN_287,
  output        _GEN_183,
  output        _GEN_256_0,
  output        _GEN_460,
  output        _GEN_278,
  output        _GEN_33,
  output        _GEN_276,
  output        _GEN_282_0,
  output        _GEN_292,
  output        _GEN_355,
  output        _GEN_48,
  output        _GEN_386,
  output        _GEN_6_1,
  output        _GEN_277_0,
  output        _GEN_21,
  output        _GEN_307,
  output        _GEN_262_0,
  output        _GEN_109,
  output        _GEN_11,
  output        _GEN_244_0,
  output        _GEN_448,
  output        _GEN_442,
  output        _GEN_21_0,
  output        _GEN_15_2,
  output        _GEN_457,
  output        _GEN_337,
  output        _GEN_30,
  output        _GEN_83,
  output        _GEN_364,
  output        _GEN_171,
  output        _GEN_186,
  output        _GEN_328,
  output        _GEN_463,
  output        _GEN_144,
  output        _GEN_279_0,
  output        _GEN_436,
  output        _GEN_97,
  output        _GEN_9_1,
  output        _GEN_264,
  output        _GEN_165,
  output        _GEN_159,
  output        _GEN_370,
  output        _GEN_250_0,
  output        _GEN_265_0,
  output        _GEN_258,
  output        _GEN_5,
  output        _GEN_285_0,
  output        _GEN_180,
  output        _GEN_271_0,
  output        _GEN_9_2,
  output        _GEN_243,
  output        _GEN_349,
  output        _GEN_343,
  output        _GEN_147,
  output        _GEN_77,
  output        _GEN_352,
  output        _GEN_174,
  output        _GEN_225,
  output        _GEN_247_0,
  output        _GEN_252,
  output        _GEN_325,
  output        _GEN_132,
  output        _GEN_147_0,
  output        _GEN_151_0,
  output        _GEN_238_0,
  output        _GEN_240,
  output        _GEN_451,
  output        _GEN_65,
  output        _GEN_273,
  output        _GEN_346,
  output        _GEN_59,
  output        _GEN_409,
  output        _GEN_231,
  output        _GEN_253_0,
  output        _GEN_331,
  output        _GEN_86,
  output        _GEN_8_0,
  output        _GEN_80,
  output        _GEN_11_0,
  output        _GEN_430,
  output        _GEN_424,
  output        _GEN_3_1,
  output        _GEN_246,
  output        _GEN_12_2,
  output        _GEN_71,
  output        _GEN_153,
  output        _GEN_168,
  output        _GEN_445,
  output        _GEN_310_0,
  output        _GEN_259_0,
  output        _GEN_267,
  output        _GEN_126,
  output        _GEN_358,
  output        _GEN_213,
  output        _GEN_255,
  output        _GEN_334,
  output        _GEN_156,
  output        _GEN_150,
  output        _GEN_412,
  output        _GEN_114,
  output        _GEN_228,
  output        _GEN_141,
  output        _GEN_11_1,
  output        _GEN_418,
  output        _GEN_427,
  output        _GEN_313_0,
  output        _GEN_292_0,
  output        _GEN_241_0,
  output        _GEN_108,
  output        _GEN_249,
  output        _GEN_6_2,
  output        _GEN_340,
  output        _GEN_312_0,
  output        _GEN_68,
  output        _GEN_74,
  output        _GEN_207,
  output        _GEN_235_0,
  output        _GEN_439,
  output        _GEN_20,
  output        _GEN_298_0,
  output        _GEN_307_0,
  output        _GEN_234,
  output        _GEN_306_0,
  output        _GEN_129,
  output        _GEN_17,
  output        _GEN_406,
  output        _GEN_89,
  output        _GEN_433,
  output        _GEN_319_0,
  output        _GEN_47,
  output        _GEN_53,
  output        _GEN_135,
  output        _GEN_391,
  output        _GEN_400,
  output        _GEN_415,
  output        _GEN_222,
  output        _GEN_295_0,
  output        _GEN_270_0,
  output        _GEN_29,
  output        _GEN_4_1,
  output        _GEN_322_0,
  output        _GEN_41,
  output        _GEN_56,
  output        _GEN_14,
  output        _GEN_195,
  output        _GEN_421,
  output        _GEN_280_0,
  output        _GEN_237,
  output        _GEN_102,
  output        _GEN_379,
  output        _GEN_62,
  output        _GEN_394,
  output        _GEN_23,
  output        _GEN_35,
  output        _GEN_123,
  output        _GEN_117,
  output        _GEN_369,
  output        _GEN_321,
  output        _GEN_216,
  output        _GEN_5_1,
  output        _GEN_14_0,
  output        _GEN_13_1,
  output        _GEN_316_0,
  output        _GEN_294_0,
  output        _GEN_50,
  output        _GEN_138,
  output        _GEN_201,
  output        _GEN_210,
  output        _GEN_96,
  output        _GEN_301_0,
  output        _GEN_315,
  output        _GEN_309,
  output        _GEN_17_0,
  output        _GEN_283_0,
  output        _GEN_273_0,
  output        _GEN_105,
  output        _GEN_382,
  output        _GEN_303,
  output        _GEN_204,
  output        _GEN_318_0,
  output        _GEN_173,
  output        _GEN_198,
  output        _GEN_258_0,
  output        _GEN_304_0,
  output        _GEN_23_0,
  output        _GEN_272_0,
  output        _GEN_120,
  output        _GEN_403,
  output        _GEN_372,
  output        _GEN_366,
  output        _GEN_267_0,
  output        _GEN_188,
  output        _GEN_289_0,
  output        _GEN_1_2,
  output        _GEN_44,
  output        _GEN_287_0,
  output        _GEN_297,
  output        _GEN_388,
  output        _GEN_397,
  output        _GEN_2_1,
  output        _GEN_252_0,
  output        _GEN_450,
  output        _GEN_99,
  output        _GEN_351,
  output        _GEN_38,
  output        _GEN_111,
  output        _GEN_219,
  output        _GEN_17_1,
  output        _GEN_7_1,
  output        _GEN_453,
  output        _GEN_447,
  output        _GEN_26,
  output        _GEN_176,
  output        _GEN_182,
  output        _GEN_438,
  output        _GEN_333,
  output        _GEN_290_0,
  output        _GEN_240_0,
  output        _GEN_0_1,
  output        _GEN_339,
  output        _GEN_32,
  output        _GEN_161,
  output        _GEN_275_0,
  output        _GEN_170,
  output        _GEN_375,
  output        _GEN_261_0,
  output        _GEN_192,
  output        _GEN_20_0,
  output        _GEN_255_0,
  output        _GEN_269_0,
  output        _GEN_10_2,
  output        _GEN_360,
  output        _GEN_281_0,
  output        _GEN_291_0,
  output        _GEN_155,
  output        _GEN_88,
  output        _GEN_300_0,
  output        _GEN_432,
  output        _GEN_11_2,
  output        _GEN_286_0,
  output        _GEN_276_0,
  output        _GEN_5_2,
  output        _GEN_254_0,
  output        _GEN_93,
  output        _GEN_5_3,
  output        _GEN_459,
  output        _GEN_385,
  output        _GEN_354,
  output        _GEN_234_0,
  output        _GEN_3_2,
  output        _GEN_146,
  output        _GEN_441,
  output        _GEN_321_0,
  output        _GEN_14_1,
  output        _GEN_257_0,
  output        _GEN_13_2,
  output        _GEN_348,
  output        _GEN_82,
  output        _GEN_357,
  output        _GEN_243_0,
  output        _GEN_8_1,
  output        _GEN_8_2,
  output        _GEN_462,
  output        _GEN_456,
  output        _GEN_342,
  output        _GEN_278_0,
  output        _GEN_70,
  output        _GEN_158,
  output        _GEN_420,
  output        _GEN_414,
  output        _GEN_236_0,
  output        _GEN_185,
  output        _GEN_336,
  output        _GEN_61,
  output        _GEN_143,
  output        _GEN_284_0,
  output        _GEN_179,
  output        _GEN_435,
  output        _GEN_242_0,
  output        _GEN_249_0,
  output        _GEN_137,
  output        _GEN_76,
  output        _GEN_164,
  output        _GEN_237_0,
  output        _GEN_315_0,
  output        _GEN_264_0,
  output        _GEN_263_0,
  output        _GEN_363,
  output        _GEN_167,
  output        _GEN_246_0,
  output        _GEN_43,
  output        _GEN_266_0,
  output        _GEN_131,
  output        _GEN_125,
  output        _GEN_317_0,
  output        _GEN_224,
  output        _GEN_150_0,
  output        _GEN_119,
  output        _GEN_239_0,
  output        _GEN_330,
  output        _GEN_152_0,
  output        _GEN_146_0,
  output        _GEN_7_2,
  output        _GEN_297_0,
  output        _GEN_245_0,
  output        _GEN_11_3,
  output        _GEN_345,
  output        _GEN_323_0,
  output        _GEN_396,
  output        _GEN_79,
  output        _GEN_218,
  output        _GEN_408,
  output        _GEN_423,
  output        _GEN_309_0,
  output        _GEN_303_0,
  output        _GEN_64,
  output        _GEN_417,
  output        _GEN_429,
  output        _GEN_444,
  output        _GEN_324,
  output        _GEN_58,
  output        _GEN_251_0,
  output        _GEN_260_0,
  output        _GEN_140,
  output        _GEN_402,
  output        _GEN_85
);
  wire  frontend_metaReset; // @[core.scala 25:25]
  wire  frontend_clock; // @[core.scala 25:25]
  wire  frontend_reset; // @[core.scala 25:25]
  wire  frontend_io_cpu_req_valid; // @[core.scala 25:25]
  wire [31:0] frontend_io_cpu_req_bits_pc; // @[core.scala 25:25]
  wire  frontend_io_cpu_resp_ready; // @[core.scala 25:25]
  wire  frontend_io_cpu_resp_valid; // @[core.scala 25:25]
  wire [31:0] frontend_io_cpu_resp_bits_pc; // @[core.scala 25:25]
  wire [31:0] frontend_io_cpu_resp_bits_inst; // @[core.scala 25:25]
  wire [31:0] frontend_io_imem_req_bits_addr; // @[core.scala 25:25]
  wire [31:0] frontend_io_imem_resp_bits_data; // @[core.scala 25:25]
  wire  frontend__GEN_1_1; // @[core.scala 25:25]
  wire  frontend__GEN_10_1; // @[core.scala 25:25]
  wire  frontend__GEN_13_1; // @[core.scala 25:25]
  wire  frontend__GEN_7_1; // @[core.scala 25:25]
  wire  frontend__GEN_9_2; // @[core.scala 25:25]
  wire  frontend__GEN_12_3; // @[core.scala 25:25]
  wire  frontend__GEN_6_3; // @[core.scala 25:25]
  wire  frontend__GEN_5_4; // @[core.scala 25:25]
  wire  frontend__GEN_8_3; // @[core.scala 25:25]
  wire  frontend__GEN_11_4; // @[core.scala 25:25]
  wire  cpath_metaReset; // @[core.scala 26:23]
  wire  cpath_clock; // @[core.scala 26:23]
  wire  cpath_io_imem_req_valid; // @[core.scala 26:23]
  wire  cpath_io_imem_resp_valid; // @[core.scala 26:23]
  wire [31:0] cpath_io_imem_resp_bits_inst; // @[core.scala 26:23]
  wire  cpath_io_dat_br_eq; // @[core.scala 26:23]
  wire  cpath_io_dat_br_lt; // @[core.scala 26:23]
  wire  cpath_io_dat_br_ltu; // @[core.scala 26:23]
  wire  cpath_io_dat_csr_eret; // @[core.scala 26:23]
  wire  cpath_io_ctl_exe_kill; // @[core.scala 26:23]
  wire [2:0] cpath_io_ctl_pc_sel; // @[core.scala 26:23]
  wire  cpath_io_ctl_brjmp_sel; // @[core.scala 26:23]
  wire [1:0] cpath_io_ctl_op1_sel; // @[core.scala 26:23]
  wire [1:0] cpath_io_ctl_op2_sel; // @[core.scala 26:23]
  wire [3:0] cpath_io_ctl_alu_fun; // @[core.scala 26:23]
  wire [1:0] cpath_io_ctl_wb_sel; // @[core.scala 26:23]
  wire  cpath_io_ctl_rf_wen; // @[core.scala 26:23]
  wire  cpath_io_ctl_bypassable; // @[core.scala 26:23]
  wire [2:0] cpath_io_ctl_csr_cmd; // @[core.scala 26:23]
  wire  cpath_io_ctl_dmem_fcn; // @[core.scala 26:23]
  wire [2:0] cpath_io_ctl_dmem_typ; // @[core.scala 26:23]
  wire  cpath_io_ctl_exception; // @[core.scala 26:23]
  wire  cpath__GEN_92_0; // @[core.scala 26:23]
  wire  cpath__GEN_52_0; // @[core.scala 26:23]
  wire  cpath__GEN_305_0; // @[core.scala 26:23]
  wire  cpath__GEN_200_0; // @[core.scala 26:23]
  wire  cpath__GEN_149_0; // @[core.scala 26:23]
  wire  cpath__GEN_25_0; // @[core.scala 26:23]
  wire  cpath__GEN_248_0; // @[core.scala 26:23]
  wire  cpath__GEN_107_0; // @[core.scala 26:23]
  wire  cpath__GEN_134_0; // @[core.scala 26:23]
  wire  cpath__GEN_206_0; // @[core.scala 26:23]
  wire  cpath__GEN_40_0; // @[core.scala 26:23]
  wire  cpath__GEN_233_0; // @[core.scala 26:23]
  wire  cpath__GEN_128_0; // @[core.scala 26:23]
  wire  cpath__GEN_191_0; // @[core.scala 26:23]
  wire  cpath__GEN_227_0; // @[core.scala 26:23]
  wire  cpath__GEN_113_0; // @[core.scala 26:23]
  wire  cpath__GEN_46_0; // @[core.scala 26:23]
  wire  cpath__GEN_299_0; // @[core.scala 26:23]
  wire  cpath__GEN_73_0; // @[core.scala 26:23]
  wire  cpath__GEN_212_0; // @[core.scala 26:23]
  wire  cpath__GEN_31_0; // @[core.scala 26:23]
  wire  cpath__GEN_311_0; // @[core.scala 26:23]
  wire  cpath__GEN_67_0; // @[core.scala 26:23]
  wire  cpath__GEN_320_0; // @[core.scala 26:23]
  wire  cpath__GEN_215_0; // @[core.scala 26:23]
  wire  cpath__GEN_221_0; // @[core.scala 26:23]
  wire  cpath__GEN_101_0; // @[core.scala 26:23]
  wire  cpath__GEN_110_0; // @[core.scala 26:23]
  wire  cpath__GEN_283_0; // @[core.scala 26:23]
  wire  cpath__GEN_314_0; // @[core.scala 26:23]
  wire  cpath__GEN_178_0; // @[core.scala 26:23]
  wire  cpath__GEN_209_0; // @[core.scala 26:23]
  wire  cpath__GEN_28_0; // @[core.scala 26:23]
  wire  cpath__GEN_277_0; // @[core.scala 26:23]
  wire  cpath__GEN_55_0; // @[core.scala 26:23]
  wire  cpath__GEN_194_0; // @[core.scala 26:23]
  wire  cpath__GEN_13_0; // @[core.scala 26:23]
  wire  cpath__GEN_49_0; // @[core.scala 26:23]
  wire  cpath__GEN_116_0; // @[core.scala 26:23]
  wire  cpath__GEN_7_0; // @[core.scala 26:23]
  wire  cpath__GEN_34_0; // @[core.scala 26:23]
  wire  cpath__GEN_122_0; // @[core.scala 26:23]
  wire  cpath__GEN_308_0; // @[core.scala 26:23]
  wire  cpath__GEN_95_0; // @[core.scala 26:23]
  wire  cpath__GEN_230_0; // @[core.scala 26:23]
  wire  cpath__GEN_293_0; // @[core.scala 26:23]
  wire  cpath__GEN_184_0; // @[core.scala 26:23]
  wire  cpath__GEN_1_2; // @[core.scala 26:23]
  wire  cpath__GEN_197_0; // @[core.scala 26:23]
  wire  cpath__GEN_187_0; // @[core.scala 26:23]
  wire  cpath__GEN_104_0; // @[core.scala 26:23]
  wire  cpath__GEN_265_0; // @[core.scala 26:23]
  wire  cpath__GEN_296_0; // @[core.scala 26:23]
  wire  cpath__GEN_160_0; // @[core.scala 26:23]
  wire  cpath__GEN_172_0; // @[core.scala 26:23]
  wire  cpath__GEN_203_0; // @[core.scala 26:23]
  wire  cpath__GEN_271_0; // @[core.scala 26:23]
  wire  cpath__GEN_37_0; // @[core.scala 26:23]
  wire  cpath__GEN_166_0; // @[core.scala 26:23]
  wire  cpath__GEN_280_0; // @[core.scala 26:23]
  wire  cpath__GEN_286_0; // @[core.scala 26:23]
  wire  cpath__GEN_22_1; // @[core.scala 26:23]
  wire  cpath__GEN_302_0; // @[core.scala 26:23]
  wire  cpath__GEN_16_2; // @[core.scala 26:23]
  wire  cpath__GEN_10_2; // @[core.scala 26:23]
  wire  cpath__GEN_259_0; // @[core.scala 26:23]
  wire  cpath__GEN_98_0; // @[core.scala 26:23]
  wire  cpath__GEN_19_1; // @[core.scala 26:23]
  wire  cpath__GEN_148_0; // @[core.scala 26:23]
  wire  cpath__GEN_87_0; // @[core.scala 26:23]
  wire  cpath__GEN_274_0; // @[core.scala 26:23]
  wire  cpath__GEN_232_0; // @[core.scala 26:23]
  wire  cpath__GEN_190_0; // @[core.scala 26:23]
  wire  cpath__GEN_154_0; // @[core.scala 26:23]
  wire  cpath__GEN_289_0; // @[core.scala 26:23]
  wire  cpath__GEN_181_0; // @[core.scala 26:23]
  wire  cpath__GEN_253_0; // @[core.scala 26:23]
  wire  cpath__GEN_72_0; // @[core.scala 26:23]
  wire  cpath__GEN_175_0; // @[core.scala 26:23]
  wire  cpath__GEN_169_0; // @[core.scala 26:23]
  wire  cpath__GEN_4_1; // @[core.scala 26:23]
  wire  cpath__GEN_247_0; // @[core.scala 26:23]
  wire  cpath__GEN_268_0; // @[core.scala 26:23]
  wire  cpath__GEN_214_0; // @[core.scala 26:23]
  wire  cpath__GEN_250_0; // @[core.scala 26:23]
  wire  cpath__GEN_241_0; // @[core.scala 26:23]
  wire  cpath__GEN_142_0; // @[core.scala 26:23]
  wire  cpath__GEN_136_0; // @[core.scala 26:23]
  wire  cpath__GEN_235_0; // @[core.scala 26:23]
  wire  cpath__GEN_262_0; // @[core.scala 26:23]
  wire  cpath__GEN_54_0; // @[core.scala 26:23]
  wire  cpath__GEN_313_0; // @[core.scala 26:23]
  wire  cpath__GEN_69_0; // @[core.scala 26:23]
  wire  cpath__GEN_157_0; // @[core.scala 26:23]
  wire  cpath__GEN_75_0; // @[core.scala 26:23]
  wire  cpath__GEN_90_0; // @[core.scala 26:23]
  wire  cpath__GEN_163_0; // @[core.scala 26:23]
  wire  cpath__GEN_130_0; // @[core.scala 26:23]
  wire  cpath__GEN_229_0; // @[core.scala 26:23]
  wire  cpath__GEN_121_0; // @[core.scala 26:23]
  wire  cpath__GEN_256_0; // @[core.scala 26:23]
  wire  cpath__GEN_81_0; // @[core.scala 26:23]
  wire  cpath__GEN_57_0; // @[core.scala 26:23]
  wire  cpath__GEN_145_0; // @[core.scala 26:23]
  wire  cpath__GEN_223_0; // @[core.scala 26:23]
  wire  cpath__GEN_118_0; // @[core.scala 26:23]
  wire  cpath__GEN_322_0; // @[core.scala 26:23]
  wire  cpath__GEN_244_0; // @[core.scala 26:23]
  wire  cpath__GEN_124_0; // @[core.scala 26:23]
  wire  cpath__GEN_103_0; // @[core.scala 26:23]
  wire  cpath__GEN_238_0; // @[core.scala 26:23]
  wire  cpath__GEN_63_0; // @[core.scala 26:23]
  wire  cpath__GEN_151_0; // @[core.scala 26:23]
  wire  cpath__GEN_202_0; // @[core.scala 26:23]
  wire  cpath__GEN_196_0; // @[core.scala 26:23]
  wire  cpath__GEN_295_0; // @[core.scala 26:23]
  wire  cpath__GEN_301_0; // @[core.scala 26:23]
  wire  cpath__GEN_310_0; // @[core.scala 26:23]
  wire  cpath__GEN_78_0; // @[core.scala 26:23]
  wire  cpath__GEN_84_0; // @[core.scala 26:23]
  wire  cpath__GEN_217_0; // @[core.scala 26:23]
  wire  cpath__GEN_36_0; // @[core.scala 26:23]
  wire  cpath__GEN_42_0; // @[core.scala 26:23]
  wire  cpath__GEN_316_0; // @[core.scala 26:23]
  wire  cpath__GEN_139_0; // @[core.scala 26:23]
  wire  cpath__GEN_18_1; // @[core.scala 26:23]
  wire  cpath__GEN_226_0; // @[core.scala 26:23]
  wire  cpath__GEN_106_0; // @[core.scala 26:23]
  wire  cpath__GEN_51_0; // @[core.scala 26:23]
  wire  cpath__GEN_45_0; // @[core.scala 26:23]
  wire  cpath__GEN_319_0; // @[core.scala 26:23]
  wire  cpath__GEN_39_0; // @[core.scala 26:23]
  wire  cpath__GEN_66_0; // @[core.scala 26:23]
  wire  cpath__GEN_24_0; // @[core.scala 26:23]
  wire  cpath__GEN_112_0; // @[core.scala 26:23]
  wire  cpath__GEN_211_0; // @[core.scala 26:23]
  wire  cpath__GEN_220_0; // @[core.scala 26:23]
  wire  cpath__GEN_133_0; // @[core.scala 26:23]
  wire  cpath__GEN_127_0; // @[core.scala 26:23]
  wire  cpath__GEN_288_1; // @[core.scala 26:23]
  wire  cpath__GEN_91_0; // @[core.scala 26:23]
  wire  cpath__GEN_205_0; // @[core.scala 26:23]
  wire  cpath__GEN_100_0; // @[core.scala 26:23]
  wire  cpath__GEN_304_0; // @[core.scala 26:23]
  wire  cpath__GEN_60_0; // @[core.scala 26:23]
  wire  cpath__GEN_298_0; // @[core.scala 26:23]
  wire  cpath__GEN_189_0; // @[core.scala 26:23]
  wire  cpath__GEN_199_0; // @[core.scala 26:23]
  wire  cpath__GEN_177_0; // @[core.scala 26:23]
  wire  cpath__GEN_12_2; // @[core.scala 26:23]
  wire  cpath__GEN_94_0; // @[core.scala 26:23]
  wire  cpath__GEN_162_0; // @[core.scala 26:23]
  wire  cpath__GEN_193_0; // @[core.scala 26:23]
  wire  cpath__GEN_208_0; // @[core.scala 26:23]
  wire  cpath__GEN_261_0; // @[core.scala 26:23]
  wire  cpath__GEN_115_0; // @[core.scala 26:23]
  wire  cpath__GEN_27_0; // @[core.scala 26:23]
  wire  cpath__GEN_270_0; // @[core.scala 26:23]
  wire  cpath__GEN_183_0; // @[core.scala 26:23]
  wire  cpath__GEN_33_0; // @[core.scala 26:23]
  wire  cpath__GEN_276_0; // @[core.scala 26:23]
  wire  cpath__GEN_282_1; // @[core.scala 26:23]
  wire  cpath__GEN_292_0; // @[core.scala 26:23]
  wire  cpath__GEN_48_0; // @[core.scala 26:23]
  wire  cpath__GEN_6_2; // @[core.scala 26:23]
  wire  cpath__GEN_307_0; // @[core.scala 26:23]
  wire  cpath__GEN_109_0; // @[core.scala 26:23]
  wire  cpath__GEN_21_1; // @[core.scala 26:23]
  wire  cpath__GEN_15_3; // @[core.scala 26:23]
  wire  cpath__GEN_30_0; // @[core.scala 26:23]
  wire  cpath__GEN_83_0; // @[core.scala 26:23]
  wire  cpath__GEN_171_0; // @[core.scala 26:23]
  wire  cpath__GEN_186_0; // @[core.scala 26:23]
  wire  cpath__GEN_144_0; // @[core.scala 26:23]
  wire  cpath__GEN_279_1; // @[core.scala 26:23]
  wire  cpath__GEN_97_0; // @[core.scala 26:23]
  wire  cpath__GEN_264_0; // @[core.scala 26:23]
  wire  cpath__GEN_165_0; // @[core.scala 26:23]
  wire  cpath__GEN_159_0; // @[core.scala 26:23]
  wire  cpath__GEN_258_0; // @[core.scala 26:23]
  wire  cpath__GEN_285_1; // @[core.scala 26:23]
  wire  cpath__GEN_180_0; // @[core.scala 26:23]
  wire  cpath__GEN_9_3; // @[core.scala 26:23]
  wire  cpath__GEN_243_0; // @[core.scala 26:23]
  wire  cpath__GEN_77_0; // @[core.scala 26:23]
  wire  cpath__GEN_174_0; // @[core.scala 26:23]
  wire  cpath__GEN_225_0; // @[core.scala 26:23]
  wire  cpath__GEN_252_0; // @[core.scala 26:23]
  wire  cpath__GEN_132_0; // @[core.scala 26:23]
  wire  cpath__GEN_147_1; // @[core.scala 26:23]
  wire  cpath__GEN_240_0; // @[core.scala 26:23]
  wire  cpath__GEN_65_0; // @[core.scala 26:23]
  wire  cpath__GEN_273_0; // @[core.scala 26:23]
  wire  cpath__GEN_59_0; // @[core.scala 26:23]
  wire  cpath__GEN_231_0; // @[core.scala 26:23]
  wire  cpath__GEN_86_0; // @[core.scala 26:23]
  wire  cpath__GEN_80_0; // @[core.scala 26:23]
  wire  cpath__GEN_3_2; // @[core.scala 26:23]
  wire  cpath__GEN_246_0; // @[core.scala 26:23]
  wire  cpath__GEN_71_0; // @[core.scala 26:23]
  wire  cpath__GEN_153_0; // @[core.scala 26:23]
  wire  cpath__GEN_168_0; // @[core.scala 26:23]
  wire  cpath__GEN_267_0; // @[core.scala 26:23]
  wire  cpath__GEN_126_0; // @[core.scala 26:23]
  wire  cpath__GEN_213_0; // @[core.scala 26:23]
  wire  cpath__GEN_255_0; // @[core.scala 26:23]
  wire  cpath__GEN_156_0; // @[core.scala 26:23]
  wire  cpath__GEN_150_0; // @[core.scala 26:23]
  wire  cpath__GEN_114_0; // @[core.scala 26:23]
  wire  cpath__GEN_228_0; // @[core.scala 26:23]
  wire  cpath__GEN_141_0; // @[core.scala 26:23]
  wire  cpath__GEN_108_0; // @[core.scala 26:23]
  wire  cpath__GEN_249_0; // @[core.scala 26:23]
  wire  cpath__GEN_312_1; // @[core.scala 26:23]
  wire  cpath__GEN_68_0; // @[core.scala 26:23]
  wire  cpath__GEN_74_0; // @[core.scala 26:23]
  wire  cpath__GEN_207_0; // @[core.scala 26:23]
  wire  cpath__GEN_234_0; // @[core.scala 26:23]
  wire  cpath__GEN_306_1; // @[core.scala 26:23]
  wire  cpath__GEN_129_0; // @[core.scala 26:23]
  wire  cpath__GEN_89_0; // @[core.scala 26:23]
  wire  cpath__GEN_47_0; // @[core.scala 26:23]
  wire  cpath__GEN_53_0; // @[core.scala 26:23]
  wire  cpath__GEN_135_0; // @[core.scala 26:23]
  wire  cpath__GEN_222_0; // @[core.scala 26:23]
  wire  cpath__GEN_29_0; // @[core.scala 26:23]
  wire  cpath__GEN_41_0; // @[core.scala 26:23]
  wire  cpath__GEN_56_0; // @[core.scala 26:23]
  wire  cpath__GEN_195_0; // @[core.scala 26:23]
  wire  cpath__GEN_237_0; // @[core.scala 26:23]
  wire  cpath__GEN_102_0; // @[core.scala 26:23]
  wire  cpath__GEN_62_0; // @[core.scala 26:23]
  wire  cpath__GEN_35_0; // @[core.scala 26:23]
  wire  cpath__GEN_123_0; // @[core.scala 26:23]
  wire  cpath__GEN_117_0; // @[core.scala 26:23]
  wire  cpath__GEN_321_0; // @[core.scala 26:23]
  wire  cpath__GEN_216_0; // @[core.scala 26:23]
  wire  cpath__GEN_294_1; // @[core.scala 26:23]
  wire  cpath__GEN_50_0; // @[core.scala 26:23]
  wire  cpath__GEN_138_0; // @[core.scala 26:23]
  wire  cpath__GEN_201_0; // @[core.scala 26:23]
  wire  cpath__GEN_210_0; // @[core.scala 26:23]
  wire  cpath__GEN_96_0; // @[core.scala 26:23]
  wire  cpath__GEN_315_0; // @[core.scala 26:23]
  wire  cpath__GEN_309_0; // @[core.scala 26:23]
  wire  cpath__GEN_17_1; // @[core.scala 26:23]
  wire  cpath__GEN_105_0; // @[core.scala 26:23]
  wire  cpath__GEN_303_0; // @[core.scala 26:23]
  wire  cpath__GEN_204_0; // @[core.scala 26:23]
  wire  cpath__GEN_318_1; // @[core.scala 26:23]
  wire  cpath__GEN_173_0; // @[core.scala 26:23]
  wire  cpath__GEN_198_0; // @[core.scala 26:23]
  wire  cpath__GEN_23_1; // @[core.scala 26:23]
  wire  cpath__GEN_272_1; // @[core.scala 26:23]
  wire  cpath__GEN_120_0; // @[core.scala 26:23]
  wire  cpath__GEN_188_0; // @[core.scala 26:23]
  wire  cpath__GEN_44_0; // @[core.scala 26:23]
  wire  cpath__GEN_287_1; // @[core.scala 26:23]
  wire  cpath__GEN_297_0; // @[core.scala 26:23]
  wire  cpath__GEN_2_2; // @[core.scala 26:23]
  wire  cpath__GEN_99_0; // @[core.scala 26:23]
  wire  cpath__GEN_38_0; // @[core.scala 26:23]
  wire  cpath__GEN_111_0; // @[core.scala 26:23]
  wire  cpath__GEN_219_0; // @[core.scala 26:23]
  wire  cpath__GEN_26_0; // @[core.scala 26:23]
  wire  cpath__GEN_176_0; // @[core.scala 26:23]
  wire  cpath__GEN_182_0; // @[core.scala 26:23]
  wire  cpath__GEN_290_1; // @[core.scala 26:23]
  wire  cpath__GEN_0_2; // @[core.scala 26:23]
  wire  cpath__GEN_32_0; // @[core.scala 26:23]
  wire  cpath__GEN_161_0; // @[core.scala 26:23]
  wire  cpath__GEN_275_1; // @[core.scala 26:23]
  wire  cpath__GEN_170_0; // @[core.scala 26:23]
  wire  cpath__GEN_192_0; // @[core.scala 26:23]
  wire  cpath__GEN_20_1; // @[core.scala 26:23]
  wire  cpath__GEN_269_1; // @[core.scala 26:23]
  wire  cpath__GEN_281_1; // @[core.scala 26:23]
  wire  cpath__GEN_291_1; // @[core.scala 26:23]
  wire  cpath__GEN_155_0; // @[core.scala 26:23]
  wire  cpath__GEN_88_0; // @[core.scala 26:23]
  wire  cpath__GEN_300_1; // @[core.scala 26:23]
  wire  cpath__GEN_11_3; // @[core.scala 26:23]
  wire  cpath__GEN_5_3; // @[core.scala 26:23]
  wire  cpath__GEN_254_1; // @[core.scala 26:23]
  wire  cpath__GEN_93_0; // @[core.scala 26:23]
  wire  cpath__GEN_14_2; // @[core.scala 26:23]
  wire  cpath__GEN_257_1; // @[core.scala 26:23]
  wire  cpath__GEN_82_0; // @[core.scala 26:23]
  wire  cpath__GEN_8_2; // @[core.scala 26:23]
  wire  cpath__GEN_278_1; // @[core.scala 26:23]
  wire  cpath__GEN_70_0; // @[core.scala 26:23]
  wire  cpath__GEN_158_0; // @[core.scala 26:23]
  wire  cpath__GEN_236_1; // @[core.scala 26:23]
  wire  cpath__GEN_185_0; // @[core.scala 26:23]
  wire  cpath__GEN_61_0; // @[core.scala 26:23]
  wire  cpath__GEN_143_0; // @[core.scala 26:23]
  wire  cpath__GEN_284_1; // @[core.scala 26:23]
  wire  cpath__GEN_179_0; // @[core.scala 26:23]
  wire  cpath__GEN_242_1; // @[core.scala 26:23]
  wire  cpath__GEN_137_0; // @[core.scala 26:23]
  wire  cpath__GEN_76_0; // @[core.scala 26:23]
  wire  cpath__GEN_164_0; // @[core.scala 26:23]
  wire  cpath__GEN_263_1; // @[core.scala 26:23]
  wire  cpath__GEN_167_0; // @[core.scala 26:23]
  wire  cpath__GEN_43_0; // @[core.scala 26:23]
  wire  cpath__GEN_266_1; // @[core.scala 26:23]
  wire  cpath__GEN_131_0; // @[core.scala 26:23]
  wire  cpath__GEN_125_0; // @[core.scala 26:23]
  wire  cpath__GEN_317_1; // @[core.scala 26:23]
  wire  cpath__GEN_224_0; // @[core.scala 26:23]
  wire  cpath__GEN_119_0; // @[core.scala 26:23]
  wire  cpath__GEN_239_1; // @[core.scala 26:23]
  wire  cpath__GEN_152_1; // @[core.scala 26:23]
  wire  cpath__GEN_146_1; // @[core.scala 26:23]
  wire  cpath__GEN_245_1; // @[core.scala 26:23]
  wire  cpath__GEN_323_1; // @[core.scala 26:23]
  wire  cpath__GEN_79_0; // @[core.scala 26:23]
  wire  cpath__GEN_218_0; // @[core.scala 26:23]
  wire  cpath__GEN_64_0; // @[core.scala 26:23]
  wire  cpath__GEN_58_0; // @[core.scala 26:23]
  wire  cpath__GEN_251_1; // @[core.scala 26:23]
  wire  cpath__GEN_260_1; // @[core.scala 26:23]
  wire  cpath__GEN_140_0; // @[core.scala 26:23]
  wire  cpath__GEN_85_0; // @[core.scala 26:23]
  wire  dpath_metaReset; // @[core.scala 27:23]
  wire  dpath_clock; // @[core.scala 27:23]
  wire  dpath_reset; // @[core.scala 27:23]
  wire [31:0] dpath_io_imem_req_bits_pc; // @[core.scala 27:23]
  wire  dpath_io_imem_resp_ready; // @[core.scala 27:23]
  wire  dpath_io_imem_resp_valid; // @[core.scala 27:23]
  wire [31:0] dpath_io_imem_resp_bits_pc; // @[core.scala 27:23]
  wire [31:0] dpath_io_imem_resp_bits_inst; // @[core.scala 27:23]
  wire [31:0] dpath_io_dmem_req_bits_addr; // @[core.scala 27:23]
  wire [31:0] dpath_io_dmem_req_bits_data; // @[core.scala 27:23]
  wire  dpath_io_dmem_req_bits_fcn; // @[core.scala 27:23]
  wire [2:0] dpath_io_dmem_req_bits_typ; // @[core.scala 27:23]
  wire [31:0] dpath_io_dmem_resp_bits_data; // @[core.scala 27:23]
  wire  dpath_io_ctl_exe_kill; // @[core.scala 27:23]
  wire [2:0] dpath_io_ctl_pc_sel; // @[core.scala 27:23]
  wire  dpath_io_ctl_brjmp_sel; // @[core.scala 27:23]
  wire [1:0] dpath_io_ctl_op1_sel; // @[core.scala 27:23]
  wire [1:0] dpath_io_ctl_op2_sel; // @[core.scala 27:23]
  wire [3:0] dpath_io_ctl_alu_fun; // @[core.scala 27:23]
  wire [1:0] dpath_io_ctl_wb_sel; // @[core.scala 27:23]
  wire  dpath_io_ctl_rf_wen; // @[core.scala 27:23]
  wire  dpath_io_ctl_bypassable; // @[core.scala 27:23]
  wire [2:0] dpath_io_ctl_csr_cmd; // @[core.scala 27:23]
  wire  dpath_io_ctl_dmem_fcn; // @[core.scala 27:23]
  wire [2:0] dpath_io_ctl_dmem_typ; // @[core.scala 27:23]
  wire  dpath_io_ctl_exception; // @[core.scala 27:23]
  wire  dpath_io_dat_br_eq; // @[core.scala 27:23]
  wire  dpath_io_dat_br_lt; // @[core.scala 27:23]
  wire  dpath_io_dat_br_ltu; // @[core.scala 27:23]
  wire  dpath_io_dat_csr_eret; // @[core.scala 27:23]
  wire  dpath__GEN_411; // @[core.scala 27:23]
  wire  dpath__GEN_405; // @[core.scala 27:23]
  wire  dpath__GEN_426; // @[core.scala 27:23]
  wire  dpath__GEN_291; // @[core.scala 27:23]
  wire  dpath__GEN_306; // @[core.scala 27:23]
  wire  dpath__GEN_384; // @[core.scala 27:23]
  wire  dpath__GEN_16_0; // @[core.scala 27:23]
  wire  dpath__GEN_19_0; // @[core.scala 27:23]
  wire  dpath__GEN_327; // @[core.scala 27:23]
  wire  dpath__GEN_390; // @[core.scala 27:23]
  wire  dpath__GEN_10_0; // @[core.scala 27:23]
  wire  dpath__GEN_285; // @[core.scala 27:23]
  wire  dpath__GEN_318; // @[core.scala 27:23]
  wire  dpath__GEN_312; // @[core.scala 27:23]
  wire  dpath__GEN_399; // @[core.scala 27:23]
  wire  dpath__GEN_387; // @[core.scala 27:23]
  wire  dpath__GEN_300; // @[core.scala 27:23]
  wire  dpath__GEN_279; // @[core.scala 27:23]
  wire  dpath__GEN_269; // @[core.scala 27:23]
  wire  dpath__GEN_378; // @[core.scala 27:23]
  wire  dpath__GEN_368; // @[core.scala 27:23]
  wire  dpath__GEN_377; // @[core.scala 27:23]
  wire  dpath__GEN_22_0; // @[core.scala 27:23]
  wire  dpath__GEN_12_0; // @[core.scala 27:23]
  wire  dpath__GEN_294; // @[core.scala 27:23]
  wire  dpath__GEN_393; // @[core.scala 27:23]
  wire  dpath__GEN_362; // @[core.scala 27:23]
  wire  dpath__GEN_461; // @[core.scala 27:23]
  wire  dpath__GEN_263; // @[core.scala 27:23]
  wire  dpath__GEN_449; // @[core.scala 27:23]
  wire  dpath__GEN_288; // @[core.scala 27:23]
  wire  dpath__GEN_245; // @[core.scala 27:23]
  wire  dpath__GEN_0_0; // @[core.scala 27:23]
  wire  dpath__GEN_272; // @[core.scala 27:23]
  wire  dpath__GEN_381; // @[core.scala 27:23]
  wire  dpath__GEN_371; // @[core.scala 27:23]
  wire  dpath__GEN_266; // @[core.scala 27:23]
  wire  dpath__GEN_16_1; // @[core.scala 27:23]
  wire  dpath__GEN_344; // @[core.scala 27:23]
  wire  dpath__GEN_282; // @[core.scala 27:23]
  wire  dpath__GEN_443; // @[core.scala 27:23]
  wire  dpath__GEN_251; // @[core.scala 27:23]
  wire  dpath__GEN_6_0; // @[core.scala 27:23]
  wire  dpath__GEN_350; // @[core.scala 27:23]
  wire  dpath__GEN_365; // @[core.scala 27:23]
  wire  dpath__GEN_15_0; // @[core.scala 27:23]
  wire  dpath__GEN_152; // @[core.scala 27:23]
  wire  dpath__GEN_446; // @[core.scala 27:23]
  wire  dpath__GEN_332; // @[core.scala 27:23]
  wire  dpath__GEN_326; // @[core.scala 27:23]
  wire  dpath__GEN_359; // @[core.scala 27:23]
  wire  dpath__GEN_15_1; // @[core.scala 27:23]
  wire  dpath__GEN_458; // @[core.scala 27:23]
  wire  dpath__GEN_452; // @[core.scala 27:23]
  wire  dpath__GEN_3_0; // @[core.scala 27:23]
  wire  dpath__GEN_347; // @[core.scala 27:23]
  wire  dpath__GEN_425; // @[core.scala 27:23]
  wire  dpath__GEN_239; // @[core.scala 27:23]
  wire  dpath__GEN_431; // @[core.scala 27:23]
  wire  dpath__GEN_254; // @[core.scala 27:23]
  wire  dpath__GEN_353; // @[core.scala 27:23]
  wire  dpath__GEN_260; // @[core.scala 27:23]
  wire  dpath__GEN_275; // @[core.scala 27:23]
  wire  dpath__GEN_9_0; // @[core.scala 27:23]
  wire  dpath__GEN_338; // @[core.scala 27:23]
  wire  dpath__GEN_374; // @[core.scala 27:23]
  wire  dpath__GEN_242; // @[core.scala 27:23]
  wire  dpath__GEN_455; // @[core.scala 27:23]
  wire  dpath__GEN_413; // @[core.scala 27:23]
  wire  dpath__GEN_236; // @[core.scala 27:23]
  wire  dpath__GEN_335; // @[core.scala 27:23]
  wire  dpath__GEN_18_0; // @[core.scala 27:23]
  wire  dpath__GEN_434; // @[core.scala 27:23]
  wire  dpath__GEN_248_0; // @[core.scala 27:23]
  wire  dpath__GEN_257; // @[core.scala 27:23]
  wire  dpath__GEN_320_0; // @[core.scala 27:23]
  wire  dpath__GEN_356; // @[core.scala 27:23]
  wire  dpath__GEN_12_1; // @[core.scala 27:23]
  wire  dpath__GEN_419; // @[core.scala 27:23]
  wire  dpath__GEN_314_0; // @[core.scala 27:23]
  wire  dpath__GEN_341; // @[core.scala 27:23]
  wire  dpath__GEN_440; // @[core.scala 27:23]
  wire  dpath__GEN_299_0; // @[core.scala 27:23]
  wire  dpath__GEN_398; // @[core.scala 27:23]
  wire  dpath__GEN_407; // @[core.scala 27:23]
  wire  dpath__GEN_149_0; // @[core.scala 27:23]
  wire  dpath__GEN_416; // @[core.scala 27:23]
  wire  dpath__GEN_281; // @[core.scala 27:23]
  wire  dpath__GEN_15_2; // @[core.scala 27:23]
  wire  dpath__GEN_380; // @[core.scala 27:23]
  wire  dpath__GEN_296_0; // @[core.scala 27:23]
  wire  dpath__GEN_422; // @[core.scala 27:23]
  wire  dpath__GEN_329; // @[core.scala 27:23]
  wire  dpath__GEN_6_1; // @[core.scala 27:23]
  wire  dpath__GEN_437; // @[core.scala 27:23]
  wire  dpath__GEN_302_0; // @[core.scala 27:23]
  wire  dpath__GEN_401; // @[core.scala 27:23]
  wire  dpath__GEN_395; // @[core.scala 27:23]
  wire  dpath__GEN_428; // @[core.scala 27:23]
  wire  dpath__GEN_308_0; // @[core.scala 27:23]
  wire  dpath__GEN_323; // @[core.scala 27:23]
  wire  dpath__GEN_317; // @[core.scala 27:23]
  wire  dpath__GEN_404; // @[core.scala 27:23]
  wire  dpath__GEN_290; // @[core.scala 27:23]
  wire  dpath__GEN_9_1; // @[core.scala 27:23]
  wire  dpath__GEN_367; // @[core.scala 27:23]
  wire  dpath__GEN_284; // @[core.scala 27:23]
  wire  dpath__GEN_274_0; // @[core.scala 27:23]
  wire  dpath__GEN_383; // @[core.scala 27:23]
  wire  dpath__GEN_373; // @[core.scala 27:23]
  wire  dpath__GEN_18_2; // @[core.scala 27:23]
  wire  dpath__GEN_410; // @[core.scala 27:23]
  wire  dpath__GEN_305_0; // @[core.scala 27:23]
  wire  dpath__GEN_8_0; // @[core.scala 27:23]
  wire  dpath__GEN_2_0; // @[core.scala 27:23]
  wire  dpath__GEN_311_0; // @[core.scala 27:23]
  wire  dpath__GEN_389; // @[core.scala 27:23]
  wire  dpath__GEN_268_0; // @[core.scala 27:23]
  wire  dpath__GEN_376; // @[core.scala 27:23]
  wire  dpath__GEN_454; // @[core.scala 27:23]
  wire  dpath__GEN_293_0; // @[core.scala 27:23]
  wire  dpath__GEN_392; // @[core.scala 27:23]
  wire  dpath__GEN_361; // @[core.scala 27:23]
  wire  dpath__GEN_287; // @[core.scala 27:23]
  wire  dpath__GEN_256_0; // @[core.scala 27:23]
  wire  dpath__GEN_460; // @[core.scala 27:23]
  wire  dpath__GEN_278; // @[core.scala 27:23]
  wire  dpath__GEN_355; // @[core.scala 27:23]
  wire  dpath__GEN_386; // @[core.scala 27:23]
  wire  dpath__GEN_277_0; // @[core.scala 27:23]
  wire  dpath__GEN_21_0; // @[core.scala 27:23]
  wire  dpath__GEN_262_0; // @[core.scala 27:23]
  wire  dpath__GEN_11_0; // @[core.scala 27:23]
  wire  dpath__GEN_244_0; // @[core.scala 27:23]
  wire  dpath__GEN_448; // @[core.scala 27:23]
  wire  dpath__GEN_442; // @[core.scala 27:23]
  wire  dpath__GEN_457; // @[core.scala 27:23]
  wire  dpath__GEN_337; // @[core.scala 27:23]
  wire  dpath__GEN_364; // @[core.scala 27:23]
  wire  dpath__GEN_328; // @[core.scala 27:23]
  wire  dpath__GEN_463; // @[core.scala 27:23]
  wire  dpath__GEN_436; // @[core.scala 27:23]
  wire  dpath__GEN_370; // @[core.scala 27:23]
  wire  dpath__GEN_250_0; // @[core.scala 27:23]
  wire  dpath__GEN_265_0; // @[core.scala 27:23]
  wire  dpath__GEN_5_0; // @[core.scala 27:23]
  wire  dpath__GEN_271_0; // @[core.scala 27:23]
  wire  dpath__GEN_349; // @[core.scala 27:23]
  wire  dpath__GEN_343; // @[core.scala 27:23]
  wire  dpath__GEN_147; // @[core.scala 27:23]
  wire  dpath__GEN_352; // @[core.scala 27:23]
  wire  dpath__GEN_247_0; // @[core.scala 27:23]
  wire  dpath__GEN_325; // @[core.scala 27:23]
  wire  dpath__GEN_151_0; // @[core.scala 27:23]
  wire  dpath__GEN_238_0; // @[core.scala 27:23]
  wire  dpath__GEN_451; // @[core.scala 27:23]
  wire  dpath__GEN_346; // @[core.scala 27:23]
  wire  dpath__GEN_409; // @[core.scala 27:23]
  wire  dpath__GEN_253_0; // @[core.scala 27:23]
  wire  dpath__GEN_331; // @[core.scala 27:23]
  wire  dpath__GEN_8_1; // @[core.scala 27:23]
  wire  dpath__GEN_11_1; // @[core.scala 27:23]
  wire  dpath__GEN_430; // @[core.scala 27:23]
  wire  dpath__GEN_424; // @[core.scala 27:23]
  wire  dpath__GEN_445; // @[core.scala 27:23]
  wire  dpath__GEN_310_0; // @[core.scala 27:23]
  wire  dpath__GEN_259_0; // @[core.scala 27:23]
  wire  dpath__GEN_358; // @[core.scala 27:23]
  wire  dpath__GEN_334; // @[core.scala 27:23]
  wire  dpath__GEN_412; // @[core.scala 27:23]
  wire  dpath__GEN_11_2; // @[core.scala 27:23]
  wire  dpath__GEN_418; // @[core.scala 27:23]
  wire  dpath__GEN_427; // @[core.scala 27:23]
  wire  dpath__GEN_313_0; // @[core.scala 27:23]
  wire  dpath__GEN_292_0; // @[core.scala 27:23]
  wire  dpath__GEN_241_0; // @[core.scala 27:23]
  wire  dpath__GEN_340; // @[core.scala 27:23]
  wire  dpath__GEN_235_0; // @[core.scala 27:23]
  wire  dpath__GEN_439; // @[core.scala 27:23]
  wire  dpath__GEN_20_0; // @[core.scala 27:23]
  wire  dpath__GEN_298_0; // @[core.scala 27:23]
  wire  dpath__GEN_307_0; // @[core.scala 27:23]
  wire  dpath__GEN_17_0; // @[core.scala 27:23]
  wire  dpath__GEN_406; // @[core.scala 27:23]
  wire  dpath__GEN_433; // @[core.scala 27:23]
  wire  dpath__GEN_319_0; // @[core.scala 27:23]
  wire  dpath__GEN_391; // @[core.scala 27:23]
  wire  dpath__GEN_400; // @[core.scala 27:23]
  wire  dpath__GEN_415; // @[core.scala 27:23]
  wire  dpath__GEN_295_0; // @[core.scala 27:23]
  wire  dpath__GEN_270_0; // @[core.scala 27:23]
  wire  dpath__GEN_4_2; // @[core.scala 27:23]
  wire  dpath__GEN_322_0; // @[core.scala 27:23]
  wire  dpath__GEN_14_0; // @[core.scala 27:23]
  wire  dpath__GEN_421; // @[core.scala 27:23]
  wire  dpath__GEN_280_0; // @[core.scala 27:23]
  wire  dpath__GEN_379; // @[core.scala 27:23]
  wire  dpath__GEN_394; // @[core.scala 27:23]
  wire  dpath__GEN_23_0; // @[core.scala 27:23]
  wire  dpath__GEN_369; // @[core.scala 27:23]
  wire  dpath__GEN_5_2; // @[core.scala 27:23]
  wire  dpath__GEN_14_1; // @[core.scala 27:23]
  wire  dpath__GEN_13_2; // @[core.scala 27:23]
  wire  dpath__GEN_316_0; // @[core.scala 27:23]
  wire  dpath__GEN_301_0; // @[core.scala 27:23]
  wire  dpath__GEN_283_0; // @[core.scala 27:23]
  wire  dpath__GEN_273_0; // @[core.scala 27:23]
  wire  dpath__GEN_382; // @[core.scala 27:23]
  wire  dpath__GEN_258_0; // @[core.scala 27:23]
  wire  dpath__GEN_304_0; // @[core.scala 27:23]
  wire  dpath__GEN_403; // @[core.scala 27:23]
  wire  dpath__GEN_372; // @[core.scala 27:23]
  wire  dpath__GEN_366; // @[core.scala 27:23]
  wire  dpath__GEN_267_0; // @[core.scala 27:23]
  wire  dpath__GEN_289_0; // @[core.scala 27:23]
  wire  dpath__GEN_1_3; // @[core.scala 27:23]
  wire  dpath__GEN_388; // @[core.scala 27:23]
  wire  dpath__GEN_397; // @[core.scala 27:23]
  wire  dpath__GEN_252_0; // @[core.scala 27:23]
  wire  dpath__GEN_450; // @[core.scala 27:23]
  wire  dpath__GEN_351; // @[core.scala 27:23]
  wire  dpath__GEN_17_2; // @[core.scala 27:23]
  wire  dpath__GEN_7_2; // @[core.scala 27:23]
  wire  dpath__GEN_453; // @[core.scala 27:23]
  wire  dpath__GEN_447; // @[core.scala 27:23]
  wire  dpath__GEN_438; // @[core.scala 27:23]
  wire  dpath__GEN_333; // @[core.scala 27:23]
  wire  dpath__GEN_240_0; // @[core.scala 27:23]
  wire  dpath__GEN_339; // @[core.scala 27:23]
  wire  dpath__GEN_375; // @[core.scala 27:23]
  wire  dpath__GEN_261_0; // @[core.scala 27:23]
  wire  dpath__GEN_255_0; // @[core.scala 27:23]
  wire  dpath__GEN_10_3; // @[core.scala 27:23]
  wire  dpath__GEN_360; // @[core.scala 27:23]
  wire  dpath__GEN_432; // @[core.scala 27:23]
  wire  dpath__GEN_286_0; // @[core.scala 27:23]
  wire  dpath__GEN_276_0; // @[core.scala 27:23]
  wire  dpath__GEN_459; // @[core.scala 27:23]
  wire  dpath__GEN_385; // @[core.scala 27:23]
  wire  dpath__GEN_354; // @[core.scala 27:23]
  wire  dpath__GEN_234_0; // @[core.scala 27:23]
  wire  dpath__GEN_3_3; // @[core.scala 27:23]
  wire  dpath__GEN_146; // @[core.scala 27:23]
  wire  dpath__GEN_441; // @[core.scala 27:23]
  wire  dpath__GEN_321_0; // @[core.scala 27:23]
  wire  dpath__GEN_13_3; // @[core.scala 27:23]
  wire  dpath__GEN_348; // @[core.scala 27:23]
  wire  dpath__GEN_357; // @[core.scala 27:23]
  wire  dpath__GEN_243_0; // @[core.scala 27:23]
  wire  dpath__GEN_462; // @[core.scala 27:23]
  wire  dpath__GEN_456; // @[core.scala 27:23]
  wire  dpath__GEN_342; // @[core.scala 27:23]
  wire  dpath__GEN_420; // @[core.scala 27:23]
  wire  dpath__GEN_414; // @[core.scala 27:23]
  wire  dpath__GEN_336; // @[core.scala 27:23]
  wire  dpath__GEN_435; // @[core.scala 27:23]
  wire  dpath__GEN_249_0; // @[core.scala 27:23]
  wire  dpath__GEN_237_0; // @[core.scala 27:23]
  wire  dpath__GEN_315_0; // @[core.scala 27:23]
  wire  dpath__GEN_264_0; // @[core.scala 27:23]
  wire  dpath__GEN_363; // @[core.scala 27:23]
  wire  dpath__GEN_246_0; // @[core.scala 27:23]
  wire  dpath__GEN_150_0; // @[core.scala 27:23]
  wire  dpath__GEN_330; // @[core.scala 27:23]
  wire  dpath__GEN_7_3; // @[core.scala 27:23]
  wire  dpath__GEN_297_0; // @[core.scala 27:23]
  wire  dpath__GEN_345; // @[core.scala 27:23]
  wire  dpath__GEN_396; // @[core.scala 27:23]
  wire  dpath__GEN_408; // @[core.scala 27:23]
  wire  dpath__GEN_423; // @[core.scala 27:23]
  wire  dpath__GEN_309_0; // @[core.scala 27:23]
  wire  dpath__GEN_303_0; // @[core.scala 27:23]
  wire  dpath__GEN_417; // @[core.scala 27:23]
  wire  dpath__GEN_429; // @[core.scala 27:23]
  wire  dpath__GEN_444; // @[core.scala 27:23]
  wire  dpath__GEN_324; // @[core.scala 27:23]
  wire  dpath__GEN_402; // @[core.scala 27:23]
  FrontEnd frontend ( // @[core.scala 25:25]
    .metaReset(frontend_metaReset),
    .clock(frontend_clock),
    .reset(frontend_reset),
    .io_cpu_req_valid(frontend_io_cpu_req_valid),
    .io_cpu_req_bits_pc(frontend_io_cpu_req_bits_pc),
    .io_cpu_resp_ready(frontend_io_cpu_resp_ready),
    .io_cpu_resp_valid(frontend_io_cpu_resp_valid),
    .io_cpu_resp_bits_pc(frontend_io_cpu_resp_bits_pc),
    .io_cpu_resp_bits_inst(frontend_io_cpu_resp_bits_inst),
    .io_imem_req_bits_addr(frontend_io_imem_req_bits_addr),
    .io_imem_resp_bits_data(frontend_io_imem_resp_bits_data),
    ._GEN_1_1(frontend__GEN_1_1),
    ._GEN_10_1(frontend__GEN_10_1),
    ._GEN_13_1(frontend__GEN_13_1),
    ._GEN_7_1(frontend__GEN_7_1),
    ._GEN_9_2(frontend__GEN_9_2),
    ._GEN_12_3(frontend__GEN_12_3),
    ._GEN_6_3(frontend__GEN_6_3),
    ._GEN_5_4(frontend__GEN_5_4),
    ._GEN_8_3(frontend__GEN_8_3),
    ._GEN_11_4(frontend__GEN_11_4)
  );
  CtlPath cpath ( // @[core.scala 26:23]
    .metaReset(cpath_metaReset),
    .clock(cpath_clock),
    .io_imem_req_valid(cpath_io_imem_req_valid),
    .io_imem_resp_valid(cpath_io_imem_resp_valid),
    .io_imem_resp_bits_inst(cpath_io_imem_resp_bits_inst),
    .io_dat_br_eq(cpath_io_dat_br_eq),
    .io_dat_br_lt(cpath_io_dat_br_lt),
    .io_dat_br_ltu(cpath_io_dat_br_ltu),
    .io_dat_csr_eret(cpath_io_dat_csr_eret),
    .io_ctl_exe_kill(cpath_io_ctl_exe_kill),
    .io_ctl_pc_sel(cpath_io_ctl_pc_sel),
    .io_ctl_brjmp_sel(cpath_io_ctl_brjmp_sel),
    .io_ctl_op1_sel(cpath_io_ctl_op1_sel),
    .io_ctl_op2_sel(cpath_io_ctl_op2_sel),
    .io_ctl_alu_fun(cpath_io_ctl_alu_fun),
    .io_ctl_wb_sel(cpath_io_ctl_wb_sel),
    .io_ctl_rf_wen(cpath_io_ctl_rf_wen),
    .io_ctl_bypassable(cpath_io_ctl_bypassable),
    .io_ctl_csr_cmd(cpath_io_ctl_csr_cmd),
    .io_ctl_dmem_fcn(cpath_io_ctl_dmem_fcn),
    .io_ctl_dmem_typ(cpath_io_ctl_dmem_typ),
    .io_ctl_exception(cpath_io_ctl_exception),
    ._GEN_92_0(cpath__GEN_92_0),
    ._GEN_52_0(cpath__GEN_52_0),
    ._GEN_305_0(cpath__GEN_305_0),
    ._GEN_200_0(cpath__GEN_200_0),
    ._GEN_149_0(cpath__GEN_149_0),
    ._GEN_25_0(cpath__GEN_25_0),
    ._GEN_248_0(cpath__GEN_248_0),
    ._GEN_107_0(cpath__GEN_107_0),
    ._GEN_134_0(cpath__GEN_134_0),
    ._GEN_206_0(cpath__GEN_206_0),
    ._GEN_40_0(cpath__GEN_40_0),
    ._GEN_233_0(cpath__GEN_233_0),
    ._GEN_128_0(cpath__GEN_128_0),
    ._GEN_191_0(cpath__GEN_191_0),
    ._GEN_227_0(cpath__GEN_227_0),
    ._GEN_113_0(cpath__GEN_113_0),
    ._GEN_46_0(cpath__GEN_46_0),
    ._GEN_299_0(cpath__GEN_299_0),
    ._GEN_73_0(cpath__GEN_73_0),
    ._GEN_212_0(cpath__GEN_212_0),
    ._GEN_31_0(cpath__GEN_31_0),
    ._GEN_311_0(cpath__GEN_311_0),
    ._GEN_67_0(cpath__GEN_67_0),
    ._GEN_320_0(cpath__GEN_320_0),
    ._GEN_215_0(cpath__GEN_215_0),
    ._GEN_221_0(cpath__GEN_221_0),
    ._GEN_101_0(cpath__GEN_101_0),
    ._GEN_110_0(cpath__GEN_110_0),
    ._GEN_283_0(cpath__GEN_283_0),
    ._GEN_314_0(cpath__GEN_314_0),
    ._GEN_178_0(cpath__GEN_178_0),
    ._GEN_209_0(cpath__GEN_209_0),
    ._GEN_28_0(cpath__GEN_28_0),
    ._GEN_277_0(cpath__GEN_277_0),
    ._GEN_55_0(cpath__GEN_55_0),
    ._GEN_194_0(cpath__GEN_194_0),
    ._GEN_13_0(cpath__GEN_13_0),
    ._GEN_49_0(cpath__GEN_49_0),
    ._GEN_116_0(cpath__GEN_116_0),
    ._GEN_7_0(cpath__GEN_7_0),
    ._GEN_34_0(cpath__GEN_34_0),
    ._GEN_122_0(cpath__GEN_122_0),
    ._GEN_308_0(cpath__GEN_308_0),
    ._GEN_95_0(cpath__GEN_95_0),
    ._GEN_230_0(cpath__GEN_230_0),
    ._GEN_293_0(cpath__GEN_293_0),
    ._GEN_184_0(cpath__GEN_184_0),
    ._GEN_1_2(cpath__GEN_1_2),
    ._GEN_197_0(cpath__GEN_197_0),
    ._GEN_187_0(cpath__GEN_187_0),
    ._GEN_104_0(cpath__GEN_104_0),
    ._GEN_265_0(cpath__GEN_265_0),
    ._GEN_296_0(cpath__GEN_296_0),
    ._GEN_160_0(cpath__GEN_160_0),
    ._GEN_172_0(cpath__GEN_172_0),
    ._GEN_203_0(cpath__GEN_203_0),
    ._GEN_271_0(cpath__GEN_271_0),
    ._GEN_37_0(cpath__GEN_37_0),
    ._GEN_166_0(cpath__GEN_166_0),
    ._GEN_280_0(cpath__GEN_280_0),
    ._GEN_286_0(cpath__GEN_286_0),
    ._GEN_22_1(cpath__GEN_22_1),
    ._GEN_302_0(cpath__GEN_302_0),
    ._GEN_16_2(cpath__GEN_16_2),
    ._GEN_10_2(cpath__GEN_10_2),
    ._GEN_259_0(cpath__GEN_259_0),
    ._GEN_98_0(cpath__GEN_98_0),
    ._GEN_19_1(cpath__GEN_19_1),
    ._GEN_148_0(cpath__GEN_148_0),
    ._GEN_87_0(cpath__GEN_87_0),
    ._GEN_274_0(cpath__GEN_274_0),
    ._GEN_232_0(cpath__GEN_232_0),
    ._GEN_190_0(cpath__GEN_190_0),
    ._GEN_154_0(cpath__GEN_154_0),
    ._GEN_289_0(cpath__GEN_289_0),
    ._GEN_181_0(cpath__GEN_181_0),
    ._GEN_253_0(cpath__GEN_253_0),
    ._GEN_72_0(cpath__GEN_72_0),
    ._GEN_175_0(cpath__GEN_175_0),
    ._GEN_169_0(cpath__GEN_169_0),
    ._GEN_4_1(cpath__GEN_4_1),
    ._GEN_247_0(cpath__GEN_247_0),
    ._GEN_268_0(cpath__GEN_268_0),
    ._GEN_214_0(cpath__GEN_214_0),
    ._GEN_250_0(cpath__GEN_250_0),
    ._GEN_241_0(cpath__GEN_241_0),
    ._GEN_142_0(cpath__GEN_142_0),
    ._GEN_136_0(cpath__GEN_136_0),
    ._GEN_235_0(cpath__GEN_235_0),
    ._GEN_262_0(cpath__GEN_262_0),
    ._GEN_54_0(cpath__GEN_54_0),
    ._GEN_313_0(cpath__GEN_313_0),
    ._GEN_69_0(cpath__GEN_69_0),
    ._GEN_157_0(cpath__GEN_157_0),
    ._GEN_75_0(cpath__GEN_75_0),
    ._GEN_90_0(cpath__GEN_90_0),
    ._GEN_163_0(cpath__GEN_163_0),
    ._GEN_130_0(cpath__GEN_130_0),
    ._GEN_229_0(cpath__GEN_229_0),
    ._GEN_121_0(cpath__GEN_121_0),
    ._GEN_256_0(cpath__GEN_256_0),
    ._GEN_81_0(cpath__GEN_81_0),
    ._GEN_57_0(cpath__GEN_57_0),
    ._GEN_145_0(cpath__GEN_145_0),
    ._GEN_223_0(cpath__GEN_223_0),
    ._GEN_118_0(cpath__GEN_118_0),
    ._GEN_322_0(cpath__GEN_322_0),
    ._GEN_244_0(cpath__GEN_244_0),
    ._GEN_124_0(cpath__GEN_124_0),
    ._GEN_103_0(cpath__GEN_103_0),
    ._GEN_238_0(cpath__GEN_238_0),
    ._GEN_63_0(cpath__GEN_63_0),
    ._GEN_151_0(cpath__GEN_151_0),
    ._GEN_202_0(cpath__GEN_202_0),
    ._GEN_196_0(cpath__GEN_196_0),
    ._GEN_295_0(cpath__GEN_295_0),
    ._GEN_301_0(cpath__GEN_301_0),
    ._GEN_310_0(cpath__GEN_310_0),
    ._GEN_78_0(cpath__GEN_78_0),
    ._GEN_84_0(cpath__GEN_84_0),
    ._GEN_217_0(cpath__GEN_217_0),
    ._GEN_36_0(cpath__GEN_36_0),
    ._GEN_42_0(cpath__GEN_42_0),
    ._GEN_316_0(cpath__GEN_316_0),
    ._GEN_139_0(cpath__GEN_139_0),
    ._GEN_18_1(cpath__GEN_18_1),
    ._GEN_226_0(cpath__GEN_226_0),
    ._GEN_106_0(cpath__GEN_106_0),
    ._GEN_51_0(cpath__GEN_51_0),
    ._GEN_45_0(cpath__GEN_45_0),
    ._GEN_319_0(cpath__GEN_319_0),
    ._GEN_39_0(cpath__GEN_39_0),
    ._GEN_66_0(cpath__GEN_66_0),
    ._GEN_24_0(cpath__GEN_24_0),
    ._GEN_112_0(cpath__GEN_112_0),
    ._GEN_211_0(cpath__GEN_211_0),
    ._GEN_220_0(cpath__GEN_220_0),
    ._GEN_133_0(cpath__GEN_133_0),
    ._GEN_127_0(cpath__GEN_127_0),
    ._GEN_288_1(cpath__GEN_288_1),
    ._GEN_91_0(cpath__GEN_91_0),
    ._GEN_205_0(cpath__GEN_205_0),
    ._GEN_100_0(cpath__GEN_100_0),
    ._GEN_304_0(cpath__GEN_304_0),
    ._GEN_60_0(cpath__GEN_60_0),
    ._GEN_298_0(cpath__GEN_298_0),
    ._GEN_189_0(cpath__GEN_189_0),
    ._GEN_199_0(cpath__GEN_199_0),
    ._GEN_177_0(cpath__GEN_177_0),
    ._GEN_12_2(cpath__GEN_12_2),
    ._GEN_94_0(cpath__GEN_94_0),
    ._GEN_162_0(cpath__GEN_162_0),
    ._GEN_193_0(cpath__GEN_193_0),
    ._GEN_208_0(cpath__GEN_208_0),
    ._GEN_261_0(cpath__GEN_261_0),
    ._GEN_115_0(cpath__GEN_115_0),
    ._GEN_27_0(cpath__GEN_27_0),
    ._GEN_270_0(cpath__GEN_270_0),
    ._GEN_183_0(cpath__GEN_183_0),
    ._GEN_33_0(cpath__GEN_33_0),
    ._GEN_276_0(cpath__GEN_276_0),
    ._GEN_282_1(cpath__GEN_282_1),
    ._GEN_292_0(cpath__GEN_292_0),
    ._GEN_48_0(cpath__GEN_48_0),
    ._GEN_6_2(cpath__GEN_6_2),
    ._GEN_307_0(cpath__GEN_307_0),
    ._GEN_109_0(cpath__GEN_109_0),
    ._GEN_21_1(cpath__GEN_21_1),
    ._GEN_15_3(cpath__GEN_15_3),
    ._GEN_30_0(cpath__GEN_30_0),
    ._GEN_83_0(cpath__GEN_83_0),
    ._GEN_171_0(cpath__GEN_171_0),
    ._GEN_186_0(cpath__GEN_186_0),
    ._GEN_144_0(cpath__GEN_144_0),
    ._GEN_279_1(cpath__GEN_279_1),
    ._GEN_97_0(cpath__GEN_97_0),
    ._GEN_264_0(cpath__GEN_264_0),
    ._GEN_165_0(cpath__GEN_165_0),
    ._GEN_159_0(cpath__GEN_159_0),
    ._GEN_258_0(cpath__GEN_258_0),
    ._GEN_285_1(cpath__GEN_285_1),
    ._GEN_180_0(cpath__GEN_180_0),
    ._GEN_9_3(cpath__GEN_9_3),
    ._GEN_243_0(cpath__GEN_243_0),
    ._GEN_77_0(cpath__GEN_77_0),
    ._GEN_174_0(cpath__GEN_174_0),
    ._GEN_225_0(cpath__GEN_225_0),
    ._GEN_252_0(cpath__GEN_252_0),
    ._GEN_132_0(cpath__GEN_132_0),
    ._GEN_147_1(cpath__GEN_147_1),
    ._GEN_240_0(cpath__GEN_240_0),
    ._GEN_65_0(cpath__GEN_65_0),
    ._GEN_273_0(cpath__GEN_273_0),
    ._GEN_59_0(cpath__GEN_59_0),
    ._GEN_231_0(cpath__GEN_231_0),
    ._GEN_86_0(cpath__GEN_86_0),
    ._GEN_80_0(cpath__GEN_80_0),
    ._GEN_3_2(cpath__GEN_3_2),
    ._GEN_246_0(cpath__GEN_246_0),
    ._GEN_71_0(cpath__GEN_71_0),
    ._GEN_153_0(cpath__GEN_153_0),
    ._GEN_168_0(cpath__GEN_168_0),
    ._GEN_267_0(cpath__GEN_267_0),
    ._GEN_126_0(cpath__GEN_126_0),
    ._GEN_213_0(cpath__GEN_213_0),
    ._GEN_255_0(cpath__GEN_255_0),
    ._GEN_156_0(cpath__GEN_156_0),
    ._GEN_150_0(cpath__GEN_150_0),
    ._GEN_114_0(cpath__GEN_114_0),
    ._GEN_228_0(cpath__GEN_228_0),
    ._GEN_141_0(cpath__GEN_141_0),
    ._GEN_108_0(cpath__GEN_108_0),
    ._GEN_249_0(cpath__GEN_249_0),
    ._GEN_312_1(cpath__GEN_312_1),
    ._GEN_68_0(cpath__GEN_68_0),
    ._GEN_74_0(cpath__GEN_74_0),
    ._GEN_207_0(cpath__GEN_207_0),
    ._GEN_234_0(cpath__GEN_234_0),
    ._GEN_306_1(cpath__GEN_306_1),
    ._GEN_129_0(cpath__GEN_129_0),
    ._GEN_89_0(cpath__GEN_89_0),
    ._GEN_47_0(cpath__GEN_47_0),
    ._GEN_53_0(cpath__GEN_53_0),
    ._GEN_135_0(cpath__GEN_135_0),
    ._GEN_222_0(cpath__GEN_222_0),
    ._GEN_29_0(cpath__GEN_29_0),
    ._GEN_41_0(cpath__GEN_41_0),
    ._GEN_56_0(cpath__GEN_56_0),
    ._GEN_195_0(cpath__GEN_195_0),
    ._GEN_237_0(cpath__GEN_237_0),
    ._GEN_102_0(cpath__GEN_102_0),
    ._GEN_62_0(cpath__GEN_62_0),
    ._GEN_35_0(cpath__GEN_35_0),
    ._GEN_123_0(cpath__GEN_123_0),
    ._GEN_117_0(cpath__GEN_117_0),
    ._GEN_321_0(cpath__GEN_321_0),
    ._GEN_216_0(cpath__GEN_216_0),
    ._GEN_294_1(cpath__GEN_294_1),
    ._GEN_50_0(cpath__GEN_50_0),
    ._GEN_138_0(cpath__GEN_138_0),
    ._GEN_201_0(cpath__GEN_201_0),
    ._GEN_210_0(cpath__GEN_210_0),
    ._GEN_96_0(cpath__GEN_96_0),
    ._GEN_315_0(cpath__GEN_315_0),
    ._GEN_309_0(cpath__GEN_309_0),
    ._GEN_17_1(cpath__GEN_17_1),
    ._GEN_105_0(cpath__GEN_105_0),
    ._GEN_303_0(cpath__GEN_303_0),
    ._GEN_204_0(cpath__GEN_204_0),
    ._GEN_318_1(cpath__GEN_318_1),
    ._GEN_173_0(cpath__GEN_173_0),
    ._GEN_198_0(cpath__GEN_198_0),
    ._GEN_23_1(cpath__GEN_23_1),
    ._GEN_272_1(cpath__GEN_272_1),
    ._GEN_120_0(cpath__GEN_120_0),
    ._GEN_188_0(cpath__GEN_188_0),
    ._GEN_44_0(cpath__GEN_44_0),
    ._GEN_287_1(cpath__GEN_287_1),
    ._GEN_297_0(cpath__GEN_297_0),
    ._GEN_2_2(cpath__GEN_2_2),
    ._GEN_99_0(cpath__GEN_99_0),
    ._GEN_38_0(cpath__GEN_38_0),
    ._GEN_111_0(cpath__GEN_111_0),
    ._GEN_219_0(cpath__GEN_219_0),
    ._GEN_26_0(cpath__GEN_26_0),
    ._GEN_176_0(cpath__GEN_176_0),
    ._GEN_182_0(cpath__GEN_182_0),
    ._GEN_290_1(cpath__GEN_290_1),
    ._GEN_0_2(cpath__GEN_0_2),
    ._GEN_32_0(cpath__GEN_32_0),
    ._GEN_161_0(cpath__GEN_161_0),
    ._GEN_275_1(cpath__GEN_275_1),
    ._GEN_170_0(cpath__GEN_170_0),
    ._GEN_192_0(cpath__GEN_192_0),
    ._GEN_20_1(cpath__GEN_20_1),
    ._GEN_269_1(cpath__GEN_269_1),
    ._GEN_281_1(cpath__GEN_281_1),
    ._GEN_291_1(cpath__GEN_291_1),
    ._GEN_155_0(cpath__GEN_155_0),
    ._GEN_88_0(cpath__GEN_88_0),
    ._GEN_300_1(cpath__GEN_300_1),
    ._GEN_11_3(cpath__GEN_11_3),
    ._GEN_5_3(cpath__GEN_5_3),
    ._GEN_254_1(cpath__GEN_254_1),
    ._GEN_93_0(cpath__GEN_93_0),
    ._GEN_14_2(cpath__GEN_14_2),
    ._GEN_257_1(cpath__GEN_257_1),
    ._GEN_82_0(cpath__GEN_82_0),
    ._GEN_8_2(cpath__GEN_8_2),
    ._GEN_278_1(cpath__GEN_278_1),
    ._GEN_70_0(cpath__GEN_70_0),
    ._GEN_158_0(cpath__GEN_158_0),
    ._GEN_236_1(cpath__GEN_236_1),
    ._GEN_185_0(cpath__GEN_185_0),
    ._GEN_61_0(cpath__GEN_61_0),
    ._GEN_143_0(cpath__GEN_143_0),
    ._GEN_284_1(cpath__GEN_284_1),
    ._GEN_179_0(cpath__GEN_179_0),
    ._GEN_242_1(cpath__GEN_242_1),
    ._GEN_137_0(cpath__GEN_137_0),
    ._GEN_76_0(cpath__GEN_76_0),
    ._GEN_164_0(cpath__GEN_164_0),
    ._GEN_263_1(cpath__GEN_263_1),
    ._GEN_167_0(cpath__GEN_167_0),
    ._GEN_43_0(cpath__GEN_43_0),
    ._GEN_266_1(cpath__GEN_266_1),
    ._GEN_131_0(cpath__GEN_131_0),
    ._GEN_125_0(cpath__GEN_125_0),
    ._GEN_317_1(cpath__GEN_317_1),
    ._GEN_224_0(cpath__GEN_224_0),
    ._GEN_119_0(cpath__GEN_119_0),
    ._GEN_239_1(cpath__GEN_239_1),
    ._GEN_152_1(cpath__GEN_152_1),
    ._GEN_146_1(cpath__GEN_146_1),
    ._GEN_245_1(cpath__GEN_245_1),
    ._GEN_323_1(cpath__GEN_323_1),
    ._GEN_79_0(cpath__GEN_79_0),
    ._GEN_218_0(cpath__GEN_218_0),
    ._GEN_64_0(cpath__GEN_64_0),
    ._GEN_58_0(cpath__GEN_58_0),
    ._GEN_251_1(cpath__GEN_251_1),
    ._GEN_260_1(cpath__GEN_260_1),
    ._GEN_140_0(cpath__GEN_140_0),
    ._GEN_85_0(cpath__GEN_85_0)
  );
  DatPath dpath ( // @[core.scala 27:23]
    .metaReset(dpath_metaReset),
    .clock(dpath_clock),
    .reset(dpath_reset),
    .io_imem_req_bits_pc(dpath_io_imem_req_bits_pc),
    .io_imem_resp_ready(dpath_io_imem_resp_ready),
    .io_imem_resp_valid(dpath_io_imem_resp_valid),
    .io_imem_resp_bits_pc(dpath_io_imem_resp_bits_pc),
    .io_imem_resp_bits_inst(dpath_io_imem_resp_bits_inst),
    .io_dmem_req_bits_addr(dpath_io_dmem_req_bits_addr),
    .io_dmem_req_bits_data(dpath_io_dmem_req_bits_data),
    .io_dmem_req_bits_fcn(dpath_io_dmem_req_bits_fcn),
    .io_dmem_req_bits_typ(dpath_io_dmem_req_bits_typ),
    .io_dmem_resp_bits_data(dpath_io_dmem_resp_bits_data),
    .io_ctl_exe_kill(dpath_io_ctl_exe_kill),
    .io_ctl_pc_sel(dpath_io_ctl_pc_sel),
    .io_ctl_brjmp_sel(dpath_io_ctl_brjmp_sel),
    .io_ctl_op1_sel(dpath_io_ctl_op1_sel),
    .io_ctl_op2_sel(dpath_io_ctl_op2_sel),
    .io_ctl_alu_fun(dpath_io_ctl_alu_fun),
    .io_ctl_wb_sel(dpath_io_ctl_wb_sel),
    .io_ctl_rf_wen(dpath_io_ctl_rf_wen),
    .io_ctl_bypassable(dpath_io_ctl_bypassable),
    .io_ctl_csr_cmd(dpath_io_ctl_csr_cmd),
    .io_ctl_dmem_fcn(dpath_io_ctl_dmem_fcn),
    .io_ctl_dmem_typ(dpath_io_ctl_dmem_typ),
    .io_ctl_exception(dpath_io_ctl_exception),
    .io_dat_br_eq(dpath_io_dat_br_eq),
    .io_dat_br_lt(dpath_io_dat_br_lt),
    .io_dat_br_ltu(dpath_io_dat_br_ltu),
    .io_dat_csr_eret(dpath_io_dat_csr_eret),
    ._GEN_411(dpath__GEN_411),
    ._GEN_405(dpath__GEN_405),
    ._GEN_426(dpath__GEN_426),
    ._GEN_291(dpath__GEN_291),
    ._GEN_306(dpath__GEN_306),
    ._GEN_384(dpath__GEN_384),
    ._GEN_16_0(dpath__GEN_16_0),
    ._GEN_19_0(dpath__GEN_19_0),
    ._GEN_327(dpath__GEN_327),
    ._GEN_390(dpath__GEN_390),
    ._GEN_10_0(dpath__GEN_10_0),
    ._GEN_285(dpath__GEN_285),
    ._GEN_318(dpath__GEN_318),
    ._GEN_312(dpath__GEN_312),
    ._GEN_399(dpath__GEN_399),
    ._GEN_387(dpath__GEN_387),
    ._GEN_300(dpath__GEN_300),
    ._GEN_279(dpath__GEN_279),
    ._GEN_269(dpath__GEN_269),
    ._GEN_378(dpath__GEN_378),
    ._GEN_368(dpath__GEN_368),
    ._GEN_377(dpath__GEN_377),
    ._GEN_22_0(dpath__GEN_22_0),
    ._GEN_12_0(dpath__GEN_12_0),
    ._GEN_294(dpath__GEN_294),
    ._GEN_393(dpath__GEN_393),
    ._GEN_362(dpath__GEN_362),
    ._GEN_461(dpath__GEN_461),
    ._GEN_263(dpath__GEN_263),
    ._GEN_449(dpath__GEN_449),
    ._GEN_288(dpath__GEN_288),
    ._GEN_245(dpath__GEN_245),
    ._GEN_0_0(dpath__GEN_0_0),
    ._GEN_272(dpath__GEN_272),
    ._GEN_381(dpath__GEN_381),
    ._GEN_371(dpath__GEN_371),
    ._GEN_266(dpath__GEN_266),
    ._GEN_16_1(dpath__GEN_16_1),
    ._GEN_344(dpath__GEN_344),
    ._GEN_282(dpath__GEN_282),
    ._GEN_443(dpath__GEN_443),
    ._GEN_251(dpath__GEN_251),
    ._GEN_6_0(dpath__GEN_6_0),
    ._GEN_350(dpath__GEN_350),
    ._GEN_365(dpath__GEN_365),
    ._GEN_15_0(dpath__GEN_15_0),
    ._GEN_152(dpath__GEN_152),
    ._GEN_446(dpath__GEN_446),
    ._GEN_332(dpath__GEN_332),
    ._GEN_326(dpath__GEN_326),
    ._GEN_359(dpath__GEN_359),
    ._GEN_15_1(dpath__GEN_15_1),
    ._GEN_458(dpath__GEN_458),
    ._GEN_452(dpath__GEN_452),
    ._GEN_3_0(dpath__GEN_3_0),
    ._GEN_347(dpath__GEN_347),
    ._GEN_425(dpath__GEN_425),
    ._GEN_239(dpath__GEN_239),
    ._GEN_431(dpath__GEN_431),
    ._GEN_254(dpath__GEN_254),
    ._GEN_353(dpath__GEN_353),
    ._GEN_260(dpath__GEN_260),
    ._GEN_275(dpath__GEN_275),
    ._GEN_9_0(dpath__GEN_9_0),
    ._GEN_338(dpath__GEN_338),
    ._GEN_374(dpath__GEN_374),
    ._GEN_242(dpath__GEN_242),
    ._GEN_455(dpath__GEN_455),
    ._GEN_413(dpath__GEN_413),
    ._GEN_236(dpath__GEN_236),
    ._GEN_335(dpath__GEN_335),
    ._GEN_18_0(dpath__GEN_18_0),
    ._GEN_434(dpath__GEN_434),
    ._GEN_248_0(dpath__GEN_248_0),
    ._GEN_257(dpath__GEN_257),
    ._GEN_320_0(dpath__GEN_320_0),
    ._GEN_356(dpath__GEN_356),
    ._GEN_12_1(dpath__GEN_12_1),
    ._GEN_419(dpath__GEN_419),
    ._GEN_314_0(dpath__GEN_314_0),
    ._GEN_341(dpath__GEN_341),
    ._GEN_440(dpath__GEN_440),
    ._GEN_299_0(dpath__GEN_299_0),
    ._GEN_398(dpath__GEN_398),
    ._GEN_407(dpath__GEN_407),
    ._GEN_149_0(dpath__GEN_149_0),
    ._GEN_416(dpath__GEN_416),
    ._GEN_281(dpath__GEN_281),
    ._GEN_15_2(dpath__GEN_15_2),
    ._GEN_380(dpath__GEN_380),
    ._GEN_296_0(dpath__GEN_296_0),
    ._GEN_422(dpath__GEN_422),
    ._GEN_329(dpath__GEN_329),
    ._GEN_6_1(dpath__GEN_6_1),
    ._GEN_437(dpath__GEN_437),
    ._GEN_302_0(dpath__GEN_302_0),
    ._GEN_401(dpath__GEN_401),
    ._GEN_395(dpath__GEN_395),
    ._GEN_428(dpath__GEN_428),
    ._GEN_308_0(dpath__GEN_308_0),
    ._GEN_323(dpath__GEN_323),
    ._GEN_317(dpath__GEN_317),
    ._GEN_404(dpath__GEN_404),
    ._GEN_290(dpath__GEN_290),
    ._GEN_9_1(dpath__GEN_9_1),
    ._GEN_367(dpath__GEN_367),
    ._GEN_284(dpath__GEN_284),
    ._GEN_274_0(dpath__GEN_274_0),
    ._GEN_383(dpath__GEN_383),
    ._GEN_373(dpath__GEN_373),
    ._GEN_18_2(dpath__GEN_18_2),
    ._GEN_410(dpath__GEN_410),
    ._GEN_305_0(dpath__GEN_305_0),
    ._GEN_8_0(dpath__GEN_8_0),
    ._GEN_2_0(dpath__GEN_2_0),
    ._GEN_311_0(dpath__GEN_311_0),
    ._GEN_389(dpath__GEN_389),
    ._GEN_268_0(dpath__GEN_268_0),
    ._GEN_376(dpath__GEN_376),
    ._GEN_454(dpath__GEN_454),
    ._GEN_293_0(dpath__GEN_293_0),
    ._GEN_392(dpath__GEN_392),
    ._GEN_361(dpath__GEN_361),
    ._GEN_287(dpath__GEN_287),
    ._GEN_256_0(dpath__GEN_256_0),
    ._GEN_460(dpath__GEN_460),
    ._GEN_278(dpath__GEN_278),
    ._GEN_355(dpath__GEN_355),
    ._GEN_386(dpath__GEN_386),
    ._GEN_277_0(dpath__GEN_277_0),
    ._GEN_21_0(dpath__GEN_21_0),
    ._GEN_262_0(dpath__GEN_262_0),
    ._GEN_11_0(dpath__GEN_11_0),
    ._GEN_244_0(dpath__GEN_244_0),
    ._GEN_448(dpath__GEN_448),
    ._GEN_442(dpath__GEN_442),
    ._GEN_457(dpath__GEN_457),
    ._GEN_337(dpath__GEN_337),
    ._GEN_364(dpath__GEN_364),
    ._GEN_328(dpath__GEN_328),
    ._GEN_463(dpath__GEN_463),
    ._GEN_436(dpath__GEN_436),
    ._GEN_370(dpath__GEN_370),
    ._GEN_250_0(dpath__GEN_250_0),
    ._GEN_265_0(dpath__GEN_265_0),
    ._GEN_5_0(dpath__GEN_5_0),
    ._GEN_271_0(dpath__GEN_271_0),
    ._GEN_349(dpath__GEN_349),
    ._GEN_343(dpath__GEN_343),
    ._GEN_147(dpath__GEN_147),
    ._GEN_352(dpath__GEN_352),
    ._GEN_247_0(dpath__GEN_247_0),
    ._GEN_325(dpath__GEN_325),
    ._GEN_151_0(dpath__GEN_151_0),
    ._GEN_238_0(dpath__GEN_238_0),
    ._GEN_451(dpath__GEN_451),
    ._GEN_346(dpath__GEN_346),
    ._GEN_409(dpath__GEN_409),
    ._GEN_253_0(dpath__GEN_253_0),
    ._GEN_331(dpath__GEN_331),
    ._GEN_8_1(dpath__GEN_8_1),
    ._GEN_11_1(dpath__GEN_11_1),
    ._GEN_430(dpath__GEN_430),
    ._GEN_424(dpath__GEN_424),
    ._GEN_445(dpath__GEN_445),
    ._GEN_310_0(dpath__GEN_310_0),
    ._GEN_259_0(dpath__GEN_259_0),
    ._GEN_358(dpath__GEN_358),
    ._GEN_334(dpath__GEN_334),
    ._GEN_412(dpath__GEN_412),
    ._GEN_11_2(dpath__GEN_11_2),
    ._GEN_418(dpath__GEN_418),
    ._GEN_427(dpath__GEN_427),
    ._GEN_313_0(dpath__GEN_313_0),
    ._GEN_292_0(dpath__GEN_292_0),
    ._GEN_241_0(dpath__GEN_241_0),
    ._GEN_340(dpath__GEN_340),
    ._GEN_235_0(dpath__GEN_235_0),
    ._GEN_439(dpath__GEN_439),
    ._GEN_20_0(dpath__GEN_20_0),
    ._GEN_298_0(dpath__GEN_298_0),
    ._GEN_307_0(dpath__GEN_307_0),
    ._GEN_17_0(dpath__GEN_17_0),
    ._GEN_406(dpath__GEN_406),
    ._GEN_433(dpath__GEN_433),
    ._GEN_319_0(dpath__GEN_319_0),
    ._GEN_391(dpath__GEN_391),
    ._GEN_400(dpath__GEN_400),
    ._GEN_415(dpath__GEN_415),
    ._GEN_295_0(dpath__GEN_295_0),
    ._GEN_270_0(dpath__GEN_270_0),
    ._GEN_4_2(dpath__GEN_4_2),
    ._GEN_322_0(dpath__GEN_322_0),
    ._GEN_14_0(dpath__GEN_14_0),
    ._GEN_421(dpath__GEN_421),
    ._GEN_280_0(dpath__GEN_280_0),
    ._GEN_379(dpath__GEN_379),
    ._GEN_394(dpath__GEN_394),
    ._GEN_23_0(dpath__GEN_23_0),
    ._GEN_369(dpath__GEN_369),
    ._GEN_5_2(dpath__GEN_5_2),
    ._GEN_14_1(dpath__GEN_14_1),
    ._GEN_13_2(dpath__GEN_13_2),
    ._GEN_316_0(dpath__GEN_316_0),
    ._GEN_301_0(dpath__GEN_301_0),
    ._GEN_283_0(dpath__GEN_283_0),
    ._GEN_273_0(dpath__GEN_273_0),
    ._GEN_382(dpath__GEN_382),
    ._GEN_258_0(dpath__GEN_258_0),
    ._GEN_304_0(dpath__GEN_304_0),
    ._GEN_403(dpath__GEN_403),
    ._GEN_372(dpath__GEN_372),
    ._GEN_366(dpath__GEN_366),
    ._GEN_267_0(dpath__GEN_267_0),
    ._GEN_289_0(dpath__GEN_289_0),
    ._GEN_1_3(dpath__GEN_1_3),
    ._GEN_388(dpath__GEN_388),
    ._GEN_397(dpath__GEN_397),
    ._GEN_252_0(dpath__GEN_252_0),
    ._GEN_450(dpath__GEN_450),
    ._GEN_351(dpath__GEN_351),
    ._GEN_17_2(dpath__GEN_17_2),
    ._GEN_7_2(dpath__GEN_7_2),
    ._GEN_453(dpath__GEN_453),
    ._GEN_447(dpath__GEN_447),
    ._GEN_438(dpath__GEN_438),
    ._GEN_333(dpath__GEN_333),
    ._GEN_240_0(dpath__GEN_240_0),
    ._GEN_339(dpath__GEN_339),
    ._GEN_375(dpath__GEN_375),
    ._GEN_261_0(dpath__GEN_261_0),
    ._GEN_255_0(dpath__GEN_255_0),
    ._GEN_10_3(dpath__GEN_10_3),
    ._GEN_360(dpath__GEN_360),
    ._GEN_432(dpath__GEN_432),
    ._GEN_286_0(dpath__GEN_286_0),
    ._GEN_276_0(dpath__GEN_276_0),
    ._GEN_459(dpath__GEN_459),
    ._GEN_385(dpath__GEN_385),
    ._GEN_354(dpath__GEN_354),
    ._GEN_234_0(dpath__GEN_234_0),
    ._GEN_3_3(dpath__GEN_3_3),
    ._GEN_146(dpath__GEN_146),
    ._GEN_441(dpath__GEN_441),
    ._GEN_321_0(dpath__GEN_321_0),
    ._GEN_13_3(dpath__GEN_13_3),
    ._GEN_348(dpath__GEN_348),
    ._GEN_357(dpath__GEN_357),
    ._GEN_243_0(dpath__GEN_243_0),
    ._GEN_462(dpath__GEN_462),
    ._GEN_456(dpath__GEN_456),
    ._GEN_342(dpath__GEN_342),
    ._GEN_420(dpath__GEN_420),
    ._GEN_414(dpath__GEN_414),
    ._GEN_336(dpath__GEN_336),
    ._GEN_435(dpath__GEN_435),
    ._GEN_249_0(dpath__GEN_249_0),
    ._GEN_237_0(dpath__GEN_237_0),
    ._GEN_315_0(dpath__GEN_315_0),
    ._GEN_264_0(dpath__GEN_264_0),
    ._GEN_363(dpath__GEN_363),
    ._GEN_246_0(dpath__GEN_246_0),
    ._GEN_150_0(dpath__GEN_150_0),
    ._GEN_330(dpath__GEN_330),
    ._GEN_7_3(dpath__GEN_7_3),
    ._GEN_297_0(dpath__GEN_297_0),
    ._GEN_345(dpath__GEN_345),
    ._GEN_396(dpath__GEN_396),
    ._GEN_408(dpath__GEN_408),
    ._GEN_423(dpath__GEN_423),
    ._GEN_309_0(dpath__GEN_309_0),
    ._GEN_303_0(dpath__GEN_303_0),
    ._GEN_417(dpath__GEN_417),
    ._GEN_429(dpath__GEN_429),
    ._GEN_444(dpath__GEN_444),
    ._GEN_324(dpath__GEN_324),
    ._GEN_402(dpath__GEN_402)
  );
  assign frontend_metaReset = metaReset;
  assign cpath_metaReset = metaReset;
  assign dpath_metaReset = metaReset;
  assign io_imem_req_bits_addr = frontend_io_imem_req_bits_addr; // @[core.scala 29:21]
  assign io_dmem_req_bits_addr = dpath_io_dmem_req_bits_addr; // @[core.scala 37:18 core.scala 38:18]
  assign io_dmem_req_bits_data = dpath_io_dmem_req_bits_data; // @[core.scala 37:18 core.scala 38:18]
  assign io_dmem_req_bits_fcn = dpath_io_dmem_req_bits_fcn; // @[core.scala 37:18 core.scala 38:18]
  assign io_dmem_req_bits_typ = dpath_io_dmem_req_bits_typ; // @[core.scala 37:18 core.scala 38:18]
  assign _GEN_411 = dpath__GEN_411;
  assign _GEN_405 = dpath__GEN_405;
  assign _GEN_92 = cpath__GEN_92_0;
  assign _GEN_52 = cpath__GEN_52_0;
  assign _GEN_305 = cpath__GEN_305_0;
  assign _GEN_200 = cpath__GEN_200_0;
  assign _GEN_149 = cpath__GEN_149_0;
  assign _GEN_426 = dpath__GEN_426;
  assign _GEN_291 = dpath__GEN_291;
  assign _GEN_1_0 = frontend__GEN_1_1;
  assign _GEN_25 = cpath__GEN_25_0;
  assign _GEN_248 = cpath__GEN_248_0;
  assign _GEN_107 = cpath__GEN_107_0;
  assign _GEN_134 = cpath__GEN_134_0;
  assign _GEN_206 = cpath__GEN_206_0;
  assign _GEN_40 = cpath__GEN_40_0;
  assign _GEN_306 = dpath__GEN_306;
  assign _GEN_233 = cpath__GEN_233_0;
  assign _GEN_128 = cpath__GEN_128_0;
  assign _GEN_384 = dpath__GEN_384;
  assign _GEN_191 = cpath__GEN_191_0;
  assign _GEN_16 = dpath__GEN_16_0;
  assign _GEN_227 = cpath__GEN_227_0;
  assign _GEN_19 = dpath__GEN_19_0;
  assign _GEN_327 = dpath__GEN_327;
  assign _GEN_113 = cpath__GEN_113_0;
  assign _GEN_46 = cpath__GEN_46_0;
  assign _GEN_299 = cpath__GEN_299_0;
  assign _GEN_390 = dpath__GEN_390;
  assign _GEN_73 = cpath__GEN_73_0;
  assign _GEN_212 = cpath__GEN_212_0;
  assign _GEN_10 = dpath__GEN_10_0;
  assign _GEN_285 = dpath__GEN_285;
  assign _GEN_318 = dpath__GEN_318;
  assign _GEN_312 = dpath__GEN_312;
  assign _GEN_31 = cpath__GEN_31_0;
  assign _GEN_311 = cpath__GEN_311_0;
  assign _GEN_67 = cpath__GEN_67_0;
  assign _GEN_320 = cpath__GEN_320_0;
  assign _GEN_399 = dpath__GEN_399;
  assign _GEN_215 = cpath__GEN_215_0;
  assign _GEN_221 = cpath__GEN_221_0;
  assign _GEN_101 = cpath__GEN_101_0;
  assign _GEN_110 = cpath__GEN_110_0;
  assign _GEN_387 = dpath__GEN_387;
  assign _GEN_283 = cpath__GEN_283_0;
  assign _GEN_314 = cpath__GEN_314_0;
  assign _GEN_178 = cpath__GEN_178_0;
  assign _GEN_209 = cpath__GEN_209_0;
  assign _GEN_300 = dpath__GEN_300;
  assign _GEN_279 = dpath__GEN_279;
  assign _GEN_269 = dpath__GEN_269;
  assign _GEN_28 = cpath__GEN_28_0;
  assign _GEN_277 = cpath__GEN_277_0;
  assign _GEN_378 = dpath__GEN_378;
  assign _GEN_368 = dpath__GEN_368;
  assign _GEN_55 = cpath__GEN_55_0;
  assign _GEN_377 = dpath__GEN_377;
  assign _GEN_194 = cpath__GEN_194_0;
  assign _GEN_22 = dpath__GEN_22_0;
  assign _GEN_12 = dpath__GEN_12_0;
  assign _GEN_294 = dpath__GEN_294;
  assign _GEN_13 = cpath__GEN_13_0;
  assign _GEN_49 = cpath__GEN_49_0;
  assign _GEN_116 = cpath__GEN_116_0;
  assign _GEN_393 = dpath__GEN_393;
  assign _GEN_362 = dpath__GEN_362;
  assign _GEN_7 = cpath__GEN_7_0;
  assign _GEN_461 = dpath__GEN_461;
  assign _GEN_34 = cpath__GEN_34_0;
  assign _GEN_122 = cpath__GEN_122_0;
  assign _GEN_308 = cpath__GEN_308_0;
  assign _GEN_263 = dpath__GEN_263;
  assign _GEN_95 = cpath__GEN_95_0;
  assign _GEN_230 = cpath__GEN_230_0;
  assign _GEN_293 = cpath__GEN_293_0;
  assign _GEN_184 = cpath__GEN_184_0;
  assign _GEN_1_1 = cpath__GEN_1_2;
  assign _GEN_10_0 = frontend__GEN_10_1;
  assign _GEN_197 = cpath__GEN_197_0;
  assign _GEN_187 = cpath__GEN_187_0;
  assign _GEN_449 = dpath__GEN_449;
  assign _GEN_288 = dpath__GEN_288;
  assign _GEN_104 = cpath__GEN_104_0;
  assign _GEN_265 = cpath__GEN_265_0;
  assign _GEN_296 = cpath__GEN_296_0;
  assign _GEN_160 = cpath__GEN_160_0;
  assign _GEN_172 = cpath__GEN_172_0;
  assign _GEN_203 = cpath__GEN_203_0;
  assign _GEN_245 = dpath__GEN_245;
  assign _GEN_0 = dpath__GEN_0_0;
  assign _GEN_272 = dpath__GEN_272;
  assign _GEN_271 = cpath__GEN_271_0;
  assign _GEN_37 = cpath__GEN_37_0;
  assign _GEN_166 = cpath__GEN_166_0;
  assign _GEN_280 = cpath__GEN_280_0;
  assign _GEN_286 = cpath__GEN_286_0;
  assign _GEN_381 = dpath__GEN_381;
  assign _GEN_371 = dpath__GEN_371;
  assign _GEN_266 = dpath__GEN_266;
  assign _GEN_16_0 = dpath__GEN_16_1;
  assign _GEN_22_0 = cpath__GEN_22_1;
  assign _GEN_302 = cpath__GEN_302_0;
  assign _GEN_344 = dpath__GEN_344;
  assign _GEN_282 = dpath__GEN_282;
  assign _GEN_443 = dpath__GEN_443;
  assign _GEN_16_1 = cpath__GEN_16_2;
  assign _GEN_251 = dpath__GEN_251;
  assign _GEN_10_1 = cpath__GEN_10_2;
  assign _GEN_259 = cpath__GEN_259_0;
  assign _GEN_98 = cpath__GEN_98_0;
  assign _GEN_6 = dpath__GEN_6_0;
  assign _GEN_350 = dpath__GEN_350;
  assign _GEN_365 = dpath__GEN_365;
  assign _GEN_15 = dpath__GEN_15_0;
  assign _GEN_152 = dpath__GEN_152;
  assign _GEN_446 = dpath__GEN_446;
  assign _GEN_332 = dpath__GEN_332;
  assign _GEN_326 = dpath__GEN_326;
  assign _GEN_19_0 = cpath__GEN_19_1;
  assign _GEN_148 = cpath__GEN_148_0;
  assign _GEN_359 = dpath__GEN_359;
  assign _GEN_15_0 = dpath__GEN_15_1;
  assign _GEN_87 = cpath__GEN_87_0;
  assign _GEN_458 = dpath__GEN_458;
  assign _GEN_452 = dpath__GEN_452;
  assign _GEN_13_0 = frontend__GEN_13_1;
  assign _GEN_3 = dpath__GEN_3_0;
  assign _GEN_347 = dpath__GEN_347;
  assign _GEN_274 = cpath__GEN_274_0;
  assign _GEN_425 = dpath__GEN_425;
  assign _GEN_239 = dpath__GEN_239;
  assign _GEN_232 = cpath__GEN_232_0;
  assign _GEN_190 = cpath__GEN_190_0;
  assign _GEN_154 = cpath__GEN_154_0;
  assign _GEN_289 = cpath__GEN_289_0;
  assign _GEN_431 = dpath__GEN_431;
  assign _GEN_181 = cpath__GEN_181_0;
  assign _GEN_253 = cpath__GEN_253_0;
  assign _GEN_254 = dpath__GEN_254;
  assign _GEN_353 = dpath__GEN_353;
  assign _GEN_72 = cpath__GEN_72_0;
  assign _GEN_175 = cpath__GEN_175_0;
  assign _GEN_169 = cpath__GEN_169_0;
  assign _GEN_260 = dpath__GEN_260;
  assign _GEN_4_0 = cpath__GEN_4_1;
  assign _GEN_275 = dpath__GEN_275;
  assign _GEN_247 = cpath__GEN_247_0;
  assign _GEN_268 = cpath__GEN_268_0;
  assign _GEN_9 = dpath__GEN_9_0;
  assign _GEN_338 = dpath__GEN_338;
  assign _GEN_374 = dpath__GEN_374;
  assign _GEN_242 = dpath__GEN_242;
  assign _GEN_214 = cpath__GEN_214_0;
  assign _GEN_250 = cpath__GEN_250_0;
  assign _GEN_455 = dpath__GEN_455;
  assign _GEN_241 = cpath__GEN_241_0;
  assign _GEN_142 = cpath__GEN_142_0;
  assign _GEN_136 = cpath__GEN_136_0;
  assign _GEN_413 = dpath__GEN_413;
  assign _GEN_235 = cpath__GEN_235_0;
  assign _GEN_236 = dpath__GEN_236;
  assign _GEN_262 = cpath__GEN_262_0;
  assign _GEN_335 = dpath__GEN_335;
  assign _GEN_54 = cpath__GEN_54_0;
  assign _GEN_313 = cpath__GEN_313_0;
  assign _GEN_18 = dpath__GEN_18_0;
  assign _GEN_69 = cpath__GEN_69_0;
  assign _GEN_157 = cpath__GEN_157_0;
  assign _GEN_434 = dpath__GEN_434;
  assign _GEN_248_0 = dpath__GEN_248_0;
  assign _GEN_257 = dpath__GEN_257;
  assign _GEN_320_0 = dpath__GEN_320_0;
  assign _GEN_75 = cpath__GEN_75_0;
  assign _GEN_356 = dpath__GEN_356;
  assign _GEN_12_0 = dpath__GEN_12_1;
  assign _GEN_90 = cpath__GEN_90_0;
  assign _GEN_163 = cpath__GEN_163_0;
  assign _GEN_419 = dpath__GEN_419;
  assign _GEN_314_0 = dpath__GEN_314_0;
  assign _GEN_7_0 = frontend__GEN_7_1;
  assign _GEN_130 = cpath__GEN_130_0;
  assign _GEN_341 = dpath__GEN_341;
  assign _GEN_440 = dpath__GEN_440;
  assign _GEN_229 = cpath__GEN_229_0;
  assign _GEN_299_0 = dpath__GEN_299_0;
  assign _GEN_121 = cpath__GEN_121_0;
  assign _GEN_256 = cpath__GEN_256_0;
  assign _GEN_398 = dpath__GEN_398;
  assign _GEN_81 = cpath__GEN_81_0;
  assign _GEN_407 = dpath__GEN_407;
  assign _GEN_149_0 = dpath__GEN_149_0;
  assign _GEN_416 = dpath__GEN_416;
  assign _GEN_281 = dpath__GEN_281;
  assign _GEN_15_1 = dpath__GEN_15_2;
  assign _GEN_380 = dpath__GEN_380;
  assign _GEN_57 = cpath__GEN_57_0;
  assign _GEN_145 = cpath__GEN_145_0;
  assign _GEN_296_0 = dpath__GEN_296_0;
  assign _GEN_223 = cpath__GEN_223_0;
  assign _GEN_118 = cpath__GEN_118_0;
  assign _GEN_322 = cpath__GEN_322_0;
  assign _GEN_422 = dpath__GEN_422;
  assign _GEN_244 = cpath__GEN_244_0;
  assign _GEN_124 = cpath__GEN_124_0;
  assign _GEN_103 = cpath__GEN_103_0;
  assign _GEN_238 = cpath__GEN_238_0;
  assign _GEN_329 = dpath__GEN_329;
  assign _GEN_63 = cpath__GEN_63_0;
  assign _GEN_151 = cpath__GEN_151_0;
  assign _GEN_202 = cpath__GEN_202_0;
  assign _GEN_6_0 = dpath__GEN_6_1;
  assign _GEN_196 = cpath__GEN_196_0;
  assign _GEN_437 = dpath__GEN_437;
  assign _GEN_302_0 = dpath__GEN_302_0;
  assign _GEN_295 = cpath__GEN_295_0;
  assign _GEN_301 = cpath__GEN_301_0;
  assign _GEN_310 = cpath__GEN_310_0;
  assign _GEN_401 = dpath__GEN_401;
  assign _GEN_395 = dpath__GEN_395;
  assign _GEN_78 = cpath__GEN_78_0;
  assign _GEN_84 = cpath__GEN_84_0;
  assign _GEN_217 = cpath__GEN_217_0;
  assign _GEN_428 = dpath__GEN_428;
  assign _GEN_308_0 = dpath__GEN_308_0;
  assign _GEN_323 = dpath__GEN_323;
  assign _GEN_36 = cpath__GEN_36_0;
  assign _GEN_42 = cpath__GEN_42_0;
  assign _GEN_317 = dpath__GEN_317;
  assign _GEN_316 = cpath__GEN_316_0;
  assign _GEN_139 = cpath__GEN_139_0;
  assign _GEN_404 = dpath__GEN_404;
  assign _GEN_290 = dpath__GEN_290;
  assign _GEN_18_0 = cpath__GEN_18_1;
  assign _GEN_226 = cpath__GEN_226_0;
  assign _GEN_106 = cpath__GEN_106_0;
  assign _GEN_51 = cpath__GEN_51_0;
  assign _GEN_45 = cpath__GEN_45_0;
  assign _GEN_9_0 = dpath__GEN_9_1;
  assign _GEN_367 = dpath__GEN_367;
  assign _GEN_319 = cpath__GEN_319_0;
  assign _GEN_284 = dpath__GEN_284;
  assign _GEN_274_0 = dpath__GEN_274_0;
  assign _GEN_39 = cpath__GEN_39_0;
  assign _GEN_383 = dpath__GEN_383;
  assign _GEN_373 = dpath__GEN_373;
  assign _GEN_66 = cpath__GEN_66_0;
  assign _GEN_18_1 = dpath__GEN_18_2;
  assign _GEN_410 = dpath__GEN_410;
  assign _GEN_24 = cpath__GEN_24_0;
  assign _GEN_305_0 = dpath__GEN_305_0;
  assign _GEN_112 = cpath__GEN_112_0;
  assign _GEN_211 = cpath__GEN_211_0;
  assign _GEN_220 = cpath__GEN_220_0;
  assign _GEN_8 = dpath__GEN_8_0;
  assign _GEN_2 = dpath__GEN_2_0;
  assign _GEN_311_0 = dpath__GEN_311_0;
  assign _GEN_133 = cpath__GEN_133_0;
  assign _GEN_127 = cpath__GEN_127_0;
  assign _GEN_288_0 = cpath__GEN_288_1;
  assign _GEN_389 = dpath__GEN_389;
  assign _GEN_91 = cpath__GEN_91_0;
  assign _GEN_205 = cpath__GEN_205_0;
  assign _GEN_100 = cpath__GEN_100_0;
  assign _GEN_304 = cpath__GEN_304_0;
  assign _GEN_60 = cpath__GEN_60_0;
  assign _GEN_298 = cpath__GEN_298_0;
  assign _GEN_189 = cpath__GEN_189_0;
  assign _GEN_199 = cpath__GEN_199_0;
  assign _GEN_177 = cpath__GEN_177_0;
  assign _GEN_12_1 = cpath__GEN_12_2;
  assign _GEN_268_0 = dpath__GEN_268_0;
  assign _GEN_94 = cpath__GEN_94_0;
  assign _GEN_376 = dpath__GEN_376;
  assign _GEN_162 = cpath__GEN_162_0;
  assign _GEN_193 = cpath__GEN_193_0;
  assign _GEN_208 = cpath__GEN_208_0;
  assign _GEN_454 = dpath__GEN_454;
  assign _GEN_293_0 = dpath__GEN_293_0;
  assign _GEN_261 = cpath__GEN_261_0;
  assign _GEN_115 = cpath__GEN_115_0;
  assign _GEN_27 = cpath__GEN_27_0;
  assign _GEN_270 = cpath__GEN_270_0;
  assign _GEN_392 = dpath__GEN_392;
  assign _GEN_361 = dpath__GEN_361;
  assign _GEN_287 = dpath__GEN_287;
  assign _GEN_183 = cpath__GEN_183_0;
  assign _GEN_256_0 = dpath__GEN_256_0;
  assign _GEN_460 = dpath__GEN_460;
  assign _GEN_278 = dpath__GEN_278;
  assign _GEN_33 = cpath__GEN_33_0;
  assign _GEN_276 = cpath__GEN_276_0;
  assign _GEN_282_0 = cpath__GEN_282_1;
  assign _GEN_292 = cpath__GEN_292_0;
  assign _GEN_355 = dpath__GEN_355;
  assign _GEN_48 = cpath__GEN_48_0;
  assign _GEN_386 = dpath__GEN_386;
  assign _GEN_6_1 = cpath__GEN_6_2;
  assign _GEN_277_0 = dpath__GEN_277_0;
  assign _GEN_21 = dpath__GEN_21_0;
  assign _GEN_307 = cpath__GEN_307_0;
  assign _GEN_262_0 = dpath__GEN_262_0;
  assign _GEN_109 = cpath__GEN_109_0;
  assign _GEN_11 = dpath__GEN_11_0;
  assign _GEN_244_0 = dpath__GEN_244_0;
  assign _GEN_448 = dpath__GEN_448;
  assign _GEN_442 = dpath__GEN_442;
  assign _GEN_21_0 = cpath__GEN_21_1;
  assign _GEN_15_2 = cpath__GEN_15_3;
  assign _GEN_457 = dpath__GEN_457;
  assign _GEN_337 = dpath__GEN_337;
  assign _GEN_30 = cpath__GEN_30_0;
  assign _GEN_83 = cpath__GEN_83_0;
  assign _GEN_364 = dpath__GEN_364;
  assign _GEN_171 = cpath__GEN_171_0;
  assign _GEN_186 = cpath__GEN_186_0;
  assign _GEN_328 = dpath__GEN_328;
  assign _GEN_463 = dpath__GEN_463;
  assign _GEN_144 = cpath__GEN_144_0;
  assign _GEN_279_0 = cpath__GEN_279_1;
  assign _GEN_436 = dpath__GEN_436;
  assign _GEN_97 = cpath__GEN_97_0;
  assign _GEN_9_1 = frontend__GEN_9_2;
  assign _GEN_264 = cpath__GEN_264_0;
  assign _GEN_165 = cpath__GEN_165_0;
  assign _GEN_159 = cpath__GEN_159_0;
  assign _GEN_370 = dpath__GEN_370;
  assign _GEN_250_0 = dpath__GEN_250_0;
  assign _GEN_265_0 = dpath__GEN_265_0;
  assign _GEN_258 = cpath__GEN_258_0;
  assign _GEN_5 = dpath__GEN_5_0;
  assign _GEN_285_0 = cpath__GEN_285_1;
  assign _GEN_180 = cpath__GEN_180_0;
  assign _GEN_271_0 = dpath__GEN_271_0;
  assign _GEN_9_2 = cpath__GEN_9_3;
  assign _GEN_243 = cpath__GEN_243_0;
  assign _GEN_349 = dpath__GEN_349;
  assign _GEN_343 = dpath__GEN_343;
  assign _GEN_147 = dpath__GEN_147;
  assign _GEN_77 = cpath__GEN_77_0;
  assign _GEN_352 = dpath__GEN_352;
  assign _GEN_174 = cpath__GEN_174_0;
  assign _GEN_225 = cpath__GEN_225_0;
  assign _GEN_247_0 = dpath__GEN_247_0;
  assign _GEN_252 = cpath__GEN_252_0;
  assign _GEN_325 = dpath__GEN_325;
  assign _GEN_132 = cpath__GEN_132_0;
  assign _GEN_147_0 = cpath__GEN_147_1;
  assign _GEN_151_0 = dpath__GEN_151_0;
  assign _GEN_238_0 = dpath__GEN_238_0;
  assign _GEN_240 = cpath__GEN_240_0;
  assign _GEN_451 = dpath__GEN_451;
  assign _GEN_65 = cpath__GEN_65_0;
  assign _GEN_273 = cpath__GEN_273_0;
  assign _GEN_346 = dpath__GEN_346;
  assign _GEN_59 = cpath__GEN_59_0;
  assign _GEN_409 = dpath__GEN_409;
  assign _GEN_231 = cpath__GEN_231_0;
  assign _GEN_253_0 = dpath__GEN_253_0;
  assign _GEN_331 = dpath__GEN_331;
  assign _GEN_86 = cpath__GEN_86_0;
  assign _GEN_8_0 = dpath__GEN_8_1;
  assign _GEN_80 = cpath__GEN_80_0;
  assign _GEN_11_0 = dpath__GEN_11_1;
  assign _GEN_430 = dpath__GEN_430;
  assign _GEN_424 = dpath__GEN_424;
  assign _GEN_3_1 = cpath__GEN_3_2;
  assign _GEN_246 = cpath__GEN_246_0;
  assign _GEN_12_2 = frontend__GEN_12_3;
  assign _GEN_71 = cpath__GEN_71_0;
  assign _GEN_153 = cpath__GEN_153_0;
  assign _GEN_168 = cpath__GEN_168_0;
  assign _GEN_445 = dpath__GEN_445;
  assign _GEN_310_0 = dpath__GEN_310_0;
  assign _GEN_259_0 = dpath__GEN_259_0;
  assign _GEN_267 = cpath__GEN_267_0;
  assign _GEN_126 = cpath__GEN_126_0;
  assign _GEN_358 = dpath__GEN_358;
  assign _GEN_213 = cpath__GEN_213_0;
  assign _GEN_255 = cpath__GEN_255_0;
  assign _GEN_334 = dpath__GEN_334;
  assign _GEN_156 = cpath__GEN_156_0;
  assign _GEN_150 = cpath__GEN_150_0;
  assign _GEN_412 = dpath__GEN_412;
  assign _GEN_114 = cpath__GEN_114_0;
  assign _GEN_228 = cpath__GEN_228_0;
  assign _GEN_141 = cpath__GEN_141_0;
  assign _GEN_11_1 = dpath__GEN_11_2;
  assign _GEN_418 = dpath__GEN_418;
  assign _GEN_427 = dpath__GEN_427;
  assign _GEN_313_0 = dpath__GEN_313_0;
  assign _GEN_292_0 = dpath__GEN_292_0;
  assign _GEN_241_0 = dpath__GEN_241_0;
  assign _GEN_108 = cpath__GEN_108_0;
  assign _GEN_249 = cpath__GEN_249_0;
  assign _GEN_6_2 = frontend__GEN_6_3;
  assign _GEN_340 = dpath__GEN_340;
  assign _GEN_312_0 = cpath__GEN_312_1;
  assign _GEN_68 = cpath__GEN_68_0;
  assign _GEN_74 = cpath__GEN_74_0;
  assign _GEN_207 = cpath__GEN_207_0;
  assign _GEN_235_0 = dpath__GEN_235_0;
  assign _GEN_439 = dpath__GEN_439;
  assign _GEN_20 = dpath__GEN_20_0;
  assign _GEN_298_0 = dpath__GEN_298_0;
  assign _GEN_307_0 = dpath__GEN_307_0;
  assign _GEN_234 = cpath__GEN_234_0;
  assign _GEN_306_0 = cpath__GEN_306_1;
  assign _GEN_129 = cpath__GEN_129_0;
  assign _GEN_17 = dpath__GEN_17_0;
  assign _GEN_406 = dpath__GEN_406;
  assign _GEN_89 = cpath__GEN_89_0;
  assign _GEN_433 = dpath__GEN_433;
  assign _GEN_319_0 = dpath__GEN_319_0;
  assign _GEN_47 = cpath__GEN_47_0;
  assign _GEN_53 = cpath__GEN_53_0;
  assign _GEN_135 = cpath__GEN_135_0;
  assign _GEN_391 = dpath__GEN_391;
  assign _GEN_400 = dpath__GEN_400;
  assign _GEN_415 = dpath__GEN_415;
  assign _GEN_222 = cpath__GEN_222_0;
  assign _GEN_295_0 = dpath__GEN_295_0;
  assign _GEN_270_0 = dpath__GEN_270_0;
  assign _GEN_29 = cpath__GEN_29_0;
  assign _GEN_4_1 = dpath__GEN_4_2;
  assign _GEN_322_0 = dpath__GEN_322_0;
  assign _GEN_41 = cpath__GEN_41_0;
  assign _GEN_56 = cpath__GEN_56_0;
  assign _GEN_14 = dpath__GEN_14_0;
  assign _GEN_195 = cpath__GEN_195_0;
  assign _GEN_421 = dpath__GEN_421;
  assign _GEN_280_0 = dpath__GEN_280_0;
  assign _GEN_237 = cpath__GEN_237_0;
  assign _GEN_102 = cpath__GEN_102_0;
  assign _GEN_379 = dpath__GEN_379;
  assign _GEN_62 = cpath__GEN_62_0;
  assign _GEN_394 = dpath__GEN_394;
  assign _GEN_23 = dpath__GEN_23_0;
  assign _GEN_35 = cpath__GEN_35_0;
  assign _GEN_123 = cpath__GEN_123_0;
  assign _GEN_117 = cpath__GEN_117_0;
  assign _GEN_369 = dpath__GEN_369;
  assign _GEN_321 = cpath__GEN_321_0;
  assign _GEN_216 = cpath__GEN_216_0;
  assign _GEN_5_1 = dpath__GEN_5_2;
  assign _GEN_14_0 = dpath__GEN_14_1;
  assign _GEN_13_1 = dpath__GEN_13_2;
  assign _GEN_316_0 = dpath__GEN_316_0;
  assign _GEN_294_0 = cpath__GEN_294_1;
  assign _GEN_50 = cpath__GEN_50_0;
  assign _GEN_138 = cpath__GEN_138_0;
  assign _GEN_201 = cpath__GEN_201_0;
  assign _GEN_210 = cpath__GEN_210_0;
  assign _GEN_96 = cpath__GEN_96_0;
  assign _GEN_301_0 = dpath__GEN_301_0;
  assign _GEN_315 = cpath__GEN_315_0;
  assign _GEN_309 = cpath__GEN_309_0;
  assign _GEN_17_0 = cpath__GEN_17_1;
  assign _GEN_283_0 = dpath__GEN_283_0;
  assign _GEN_273_0 = dpath__GEN_273_0;
  assign _GEN_105 = cpath__GEN_105_0;
  assign _GEN_382 = dpath__GEN_382;
  assign _GEN_303 = cpath__GEN_303_0;
  assign _GEN_204 = cpath__GEN_204_0;
  assign _GEN_318_0 = cpath__GEN_318_1;
  assign _GEN_173 = cpath__GEN_173_0;
  assign _GEN_198 = cpath__GEN_198_0;
  assign _GEN_258_0 = dpath__GEN_258_0;
  assign _GEN_304_0 = dpath__GEN_304_0;
  assign _GEN_23_0 = cpath__GEN_23_1;
  assign _GEN_272_0 = cpath__GEN_272_1;
  assign _GEN_120 = cpath__GEN_120_0;
  assign _GEN_403 = dpath__GEN_403;
  assign _GEN_372 = dpath__GEN_372;
  assign _GEN_366 = dpath__GEN_366;
  assign _GEN_267_0 = dpath__GEN_267_0;
  assign _GEN_188 = cpath__GEN_188_0;
  assign _GEN_289_0 = dpath__GEN_289_0;
  assign _GEN_1_2 = dpath__GEN_1_3;
  assign _GEN_44 = cpath__GEN_44_0;
  assign _GEN_287_0 = cpath__GEN_287_1;
  assign _GEN_297 = cpath__GEN_297_0;
  assign _GEN_388 = dpath__GEN_388;
  assign _GEN_397 = dpath__GEN_397;
  assign _GEN_2_1 = cpath__GEN_2_2;
  assign _GEN_252_0 = dpath__GEN_252_0;
  assign _GEN_450 = dpath__GEN_450;
  assign _GEN_99 = cpath__GEN_99_0;
  assign _GEN_351 = dpath__GEN_351;
  assign _GEN_38 = cpath__GEN_38_0;
  assign _GEN_111 = cpath__GEN_111_0;
  assign _GEN_219 = cpath__GEN_219_0;
  assign _GEN_17_1 = dpath__GEN_17_2;
  assign _GEN_7_1 = dpath__GEN_7_2;
  assign _GEN_453 = dpath__GEN_453;
  assign _GEN_447 = dpath__GEN_447;
  assign _GEN_26 = cpath__GEN_26_0;
  assign _GEN_176 = cpath__GEN_176_0;
  assign _GEN_182 = cpath__GEN_182_0;
  assign _GEN_438 = dpath__GEN_438;
  assign _GEN_333 = dpath__GEN_333;
  assign _GEN_290_0 = cpath__GEN_290_1;
  assign _GEN_240_0 = dpath__GEN_240_0;
  assign _GEN_0_1 = cpath__GEN_0_2;
  assign _GEN_339 = dpath__GEN_339;
  assign _GEN_32 = cpath__GEN_32_0;
  assign _GEN_161 = cpath__GEN_161_0;
  assign _GEN_275_0 = cpath__GEN_275_1;
  assign _GEN_170 = cpath__GEN_170_0;
  assign _GEN_375 = dpath__GEN_375;
  assign _GEN_261_0 = dpath__GEN_261_0;
  assign _GEN_192 = cpath__GEN_192_0;
  assign _GEN_20_0 = cpath__GEN_20_1;
  assign _GEN_255_0 = dpath__GEN_255_0;
  assign _GEN_269_0 = cpath__GEN_269_1;
  assign _GEN_10_2 = dpath__GEN_10_3;
  assign _GEN_360 = dpath__GEN_360;
  assign _GEN_281_0 = cpath__GEN_281_1;
  assign _GEN_291_0 = cpath__GEN_291_1;
  assign _GEN_155 = cpath__GEN_155_0;
  assign _GEN_88 = cpath__GEN_88_0;
  assign _GEN_300_0 = cpath__GEN_300_1;
  assign _GEN_432 = dpath__GEN_432;
  assign _GEN_11_2 = cpath__GEN_11_3;
  assign _GEN_286_0 = dpath__GEN_286_0;
  assign _GEN_276_0 = dpath__GEN_276_0;
  assign _GEN_5_2 = cpath__GEN_5_3;
  assign _GEN_254_0 = cpath__GEN_254_1;
  assign _GEN_93 = cpath__GEN_93_0;
  assign _GEN_5_3 = frontend__GEN_5_4;
  assign _GEN_459 = dpath__GEN_459;
  assign _GEN_385 = dpath__GEN_385;
  assign _GEN_354 = dpath__GEN_354;
  assign _GEN_234_0 = dpath__GEN_234_0;
  assign _GEN_3_2 = dpath__GEN_3_3;
  assign _GEN_146 = dpath__GEN_146;
  assign _GEN_441 = dpath__GEN_441;
  assign _GEN_321_0 = dpath__GEN_321_0;
  assign _GEN_14_1 = cpath__GEN_14_2;
  assign _GEN_257_0 = cpath__GEN_257_1;
  assign _GEN_13_2 = dpath__GEN_13_3;
  assign _GEN_348 = dpath__GEN_348;
  assign _GEN_82 = cpath__GEN_82_0;
  assign _GEN_357 = dpath__GEN_357;
  assign _GEN_243_0 = dpath__GEN_243_0;
  assign _GEN_8_1 = cpath__GEN_8_2;
  assign _GEN_8_2 = frontend__GEN_8_3;
  assign _GEN_462 = dpath__GEN_462;
  assign _GEN_456 = dpath__GEN_456;
  assign _GEN_342 = dpath__GEN_342;
  assign _GEN_278_0 = cpath__GEN_278_1;
  assign _GEN_70 = cpath__GEN_70_0;
  assign _GEN_158 = cpath__GEN_158_0;
  assign _GEN_420 = dpath__GEN_420;
  assign _GEN_414 = dpath__GEN_414;
  assign _GEN_236_0 = cpath__GEN_236_1;
  assign _GEN_185 = cpath__GEN_185_0;
  assign _GEN_336 = dpath__GEN_336;
  assign _GEN_61 = cpath__GEN_61_0;
  assign _GEN_143 = cpath__GEN_143_0;
  assign _GEN_284_0 = cpath__GEN_284_1;
  assign _GEN_179 = cpath__GEN_179_0;
  assign _GEN_435 = dpath__GEN_435;
  assign _GEN_242_0 = cpath__GEN_242_1;
  assign _GEN_249_0 = dpath__GEN_249_0;
  assign _GEN_137 = cpath__GEN_137_0;
  assign _GEN_76 = cpath__GEN_76_0;
  assign _GEN_164 = cpath__GEN_164_0;
  assign _GEN_237_0 = dpath__GEN_237_0;
  assign _GEN_315_0 = dpath__GEN_315_0;
  assign _GEN_264_0 = dpath__GEN_264_0;
  assign _GEN_263_0 = cpath__GEN_263_1;
  assign _GEN_363 = dpath__GEN_363;
  assign _GEN_167 = cpath__GEN_167_0;
  assign _GEN_246_0 = dpath__GEN_246_0;
  assign _GEN_43 = cpath__GEN_43_0;
  assign _GEN_266_0 = cpath__GEN_266_1;
  assign _GEN_131 = cpath__GEN_131_0;
  assign _GEN_125 = cpath__GEN_125_0;
  assign _GEN_317_0 = cpath__GEN_317_1;
  assign _GEN_224 = cpath__GEN_224_0;
  assign _GEN_150_0 = dpath__GEN_150_0;
  assign _GEN_119 = cpath__GEN_119_0;
  assign _GEN_239_0 = cpath__GEN_239_1;
  assign _GEN_330 = dpath__GEN_330;
  assign _GEN_152_0 = cpath__GEN_152_1;
  assign _GEN_146_0 = cpath__GEN_146_1;
  assign _GEN_7_2 = dpath__GEN_7_3;
  assign _GEN_297_0 = dpath__GEN_297_0;
  assign _GEN_245_0 = cpath__GEN_245_1;
  assign _GEN_11_3 = frontend__GEN_11_4;
  assign _GEN_345 = dpath__GEN_345;
  assign _GEN_323_0 = cpath__GEN_323_1;
  assign _GEN_396 = dpath__GEN_396;
  assign _GEN_79 = cpath__GEN_79_0;
  assign _GEN_218 = cpath__GEN_218_0;
  assign _GEN_408 = dpath__GEN_408;
  assign _GEN_423 = dpath__GEN_423;
  assign _GEN_309_0 = dpath__GEN_309_0;
  assign _GEN_303_0 = dpath__GEN_303_0;
  assign _GEN_64 = cpath__GEN_64_0;
  assign _GEN_417 = dpath__GEN_417;
  assign _GEN_429 = dpath__GEN_429;
  assign _GEN_444 = dpath__GEN_444;
  assign _GEN_324 = dpath__GEN_324;
  assign _GEN_58 = cpath__GEN_58_0;
  assign _GEN_251_0 = cpath__GEN_251_1;
  assign _GEN_260_0 = cpath__GEN_260_1;
  assign _GEN_140 = cpath__GEN_140_0;
  assign _GEN_402 = dpath__GEN_402;
  assign _GEN_85 = cpath__GEN_85_0;
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_io_cpu_req_valid = cpath_io_imem_req_valid; // @[core.scala 30:20 core.scala 31:20 core.scala 32:30]
  assign frontend_io_cpu_req_bits_pc = dpath_io_imem_req_bits_pc; // @[core.scala 30:20 core.scala 31:20]
  assign frontend_io_cpu_resp_ready = dpath_io_imem_resp_ready; // @[core.scala 30:20 core.scala 31:20]
  assign frontend_io_imem_resp_bits_data = io_imem_resp_bits_data; // @[core.scala 29:21]
  assign cpath_clock = clock;
  assign cpath_io_imem_resp_valid = frontend_io_cpu_resp_valid; // @[core.scala 30:20]
  assign cpath_io_imem_resp_bits_inst = frontend_io_cpu_resp_bits_inst; // @[core.scala 30:20]
  assign cpath_io_dat_br_eq = dpath_io_dat_br_eq; // @[core.scala 35:18]
  assign cpath_io_dat_br_lt = dpath_io_dat_br_lt; // @[core.scala 35:18]
  assign cpath_io_dat_br_ltu = dpath_io_dat_br_ltu; // @[core.scala 35:18]
  assign cpath_io_dat_csr_eret = dpath_io_dat_csr_eret; // @[core.scala 35:18]
  assign dpath_clock = clock;
  assign dpath_reset = reset;
  assign dpath_io_imem_resp_valid = frontend_io_cpu_resp_valid; // @[core.scala 31:20]
  assign dpath_io_imem_resp_bits_pc = frontend_io_cpu_resp_bits_pc; // @[core.scala 31:20]
  assign dpath_io_imem_resp_bits_inst = frontend_io_cpu_resp_bits_inst; // @[core.scala 31:20]
  assign dpath_io_dmem_resp_bits_data = io_dmem_resp_bits_data; // @[core.scala 38:18]
  assign dpath_io_ctl_exe_kill = cpath_io_ctl_exe_kill; // @[core.scala 34:18]
  assign dpath_io_ctl_pc_sel = cpath_io_ctl_pc_sel; // @[core.scala 34:18]
  assign dpath_io_ctl_brjmp_sel = cpath_io_ctl_brjmp_sel; // @[core.scala 34:18]
  assign dpath_io_ctl_op1_sel = cpath_io_ctl_op1_sel; // @[core.scala 34:18]
  assign dpath_io_ctl_op2_sel = cpath_io_ctl_op2_sel; // @[core.scala 34:18]
  assign dpath_io_ctl_alu_fun = cpath_io_ctl_alu_fun; // @[core.scala 34:18]
  assign dpath_io_ctl_wb_sel = cpath_io_ctl_wb_sel; // @[core.scala 34:18]
  assign dpath_io_ctl_rf_wen = cpath_io_ctl_rf_wen; // @[core.scala 34:18]
  assign dpath_io_ctl_bypassable = cpath_io_ctl_bypassable; // @[core.scala 34:18]
  assign dpath_io_ctl_csr_cmd = cpath_io_ctl_csr_cmd; // @[core.scala 34:18]
  assign dpath_io_ctl_dmem_fcn = cpath_io_ctl_dmem_fcn; // @[core.scala 34:18]
  assign dpath_io_ctl_dmem_typ = cpath_io_ctl_dmem_typ; // @[core.scala 34:18]
  assign dpath_io_ctl_exception = cpath_io_ctl_exception; // @[core.scala 34:18]
endmodule
module SyncMem(
  input         metaReset,
  input         clock,
  input  [20:0] io_dataInstr_0_addr,
  output [31:0] io_dataInstr_0_data,
  input  [20:0] io_dw_addr,
  input  [31:0] io_dw_data,
  input         io_dw_en
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  mem_sparse_metaReset; // @[memory.scala 97:36]
  wire  mem_sparse_clock; // @[memory.scala 97:36]
  wire [20:0] mem_sparse_io_w_1_addr; // @[memory.scala 97:36]
  wire  mem_sparse_io_w_1_en; // @[memory.scala 97:36]
  wire [7:0] mem_sparse_io_w_1_data; // @[memory.scala 97:36]
  wire [20:0] mem_sparse_io_r_0_addr; // @[memory.scala 97:36]
  wire [7:0] mem_sparse_io_r_0_data; // @[memory.scala 97:36]
  wire  mem_sparse_0_metaReset; // @[memory.scala 97:36]
  wire  mem_sparse_0_clock; // @[memory.scala 97:36]
  wire [20:0] mem_sparse_0_io_w_1_addr; // @[memory.scala 97:36]
  wire  mem_sparse_0_io_w_1_en; // @[memory.scala 97:36]
  wire [7:0] mem_sparse_0_io_w_1_data; // @[memory.scala 97:36]
  wire [20:0] mem_sparse_0_io_r_0_addr; // @[memory.scala 97:36]
  wire [7:0] mem_sparse_0_io_r_0_data; // @[memory.scala 97:36]
  wire  mem_sparse_1_metaReset; // @[memory.scala 97:36]
  wire  mem_sparse_1_clock; // @[memory.scala 97:36]
  wire [20:0] mem_sparse_1_io_w_1_addr; // @[memory.scala 97:36]
  wire  mem_sparse_1_io_w_1_en; // @[memory.scala 97:36]
  wire [7:0] mem_sparse_1_io_w_1_data; // @[memory.scala 97:36]
  wire [20:0] mem_sparse_1_io_r_0_addr; // @[memory.scala 97:36]
  wire [7:0] mem_sparse_1_io_r_0_data; // @[memory.scala 97:36]
  wire  mem_sparse_2_metaReset; // @[memory.scala 97:36]
  wire  mem_sparse_2_clock; // @[memory.scala 97:36]
  wire [20:0] mem_sparse_2_io_w_1_addr; // @[memory.scala 97:36]
  wire  mem_sparse_2_io_w_1_en; // @[memory.scala 97:36]
  wire [7:0] mem_sparse_2_io_w_1_data; // @[memory.scala 97:36]
  wire [20:0] mem_sparse_2_io_r_0_addr; // @[memory.scala 97:36]
  wire [7:0] mem_sparse_2_io_r_0_data; // @[memory.scala 97:36]
  reg [20:0] underlying_0__T_54_addr_pipe_0;
  reg [20:0] underlying_1__T_54_addr_pipe_0;
  reg [20:0] underlying_2__T_54_addr_pipe_0;
  reg [20:0] underlying_3__T_54_addr_pipe_0;
  wire [7:0] underlying_1__T_54_data = mem_sparse_0_io_r_0_data; // @[memory.scala 97:36]
  wire [7:0] underlying_0__T_54_data = mem_sparse_io_r_0_data; // @[memory.scala 97:36]
  wire [15:0] _T_68 = {underlying_1__T_54_data,underlying_0__T_54_data}; // @[memory.scala 82:55]
  wire [7:0] underlying_3__T_54_data = mem_sparse_2_io_r_0_data; // @[memory.scala 97:36]
  wire [7:0] underlying_2__T_54_data = mem_sparse_1_io_r_0_data; // @[memory.scala 97:36]
  wire [15:0] _T_69 = {underlying_3__T_54_data,underlying_2__T_54_data}; // @[memory.scala 82:55]
  SparseMem_0 mem_sparse ( // @[memory.scala 97:36]
    .metaReset(mem_sparse_metaReset),
    .clock(mem_sparse_clock),
    .io_w_1_addr(mem_sparse_io_w_1_addr),
    .io_w_1_en(mem_sparse_io_w_1_en),
    .io_w_1_data(mem_sparse_io_w_1_data),
    .io_r_0_addr(mem_sparse_io_r_0_addr),
    .io_r_0_data(mem_sparse_io_r_0_data)
  );
  SparseMem_0 mem_sparse_0 ( // @[memory.scala 97:36]
    .metaReset(mem_sparse_0_metaReset),
    .clock(mem_sparse_0_clock),
    .io_w_1_addr(mem_sparse_0_io_w_1_addr),
    .io_w_1_en(mem_sparse_0_io_w_1_en),
    .io_w_1_data(mem_sparse_0_io_w_1_data),
    .io_r_0_addr(mem_sparse_0_io_r_0_addr),
    .io_r_0_data(mem_sparse_0_io_r_0_data)
  );
  SparseMem_0 mem_sparse_1 ( // @[memory.scala 97:36]
    .metaReset(mem_sparse_1_metaReset),
    .clock(mem_sparse_1_clock),
    .io_w_1_addr(mem_sparse_1_io_w_1_addr),
    .io_w_1_en(mem_sparse_1_io_w_1_en),
    .io_w_1_data(mem_sparse_1_io_w_1_data),
    .io_r_0_addr(mem_sparse_1_io_r_0_addr),
    .io_r_0_data(mem_sparse_1_io_r_0_data)
  );
  SparseMem_0 mem_sparse_2 ( // @[memory.scala 97:36]
    .metaReset(mem_sparse_2_metaReset),
    .clock(mem_sparse_2_clock),
    .io_w_1_addr(mem_sparse_2_io_w_1_addr),
    .io_w_1_en(mem_sparse_2_io_w_1_en),
    .io_w_1_data(mem_sparse_2_io_w_1_data),
    .io_r_0_addr(mem_sparse_2_io_r_0_addr),
    .io_r_0_data(mem_sparse_2_io_r_0_data)
  );
  assign mem_sparse_metaReset = metaReset;
  assign mem_sparse_0_metaReset = metaReset;
  assign mem_sparse_1_metaReset = metaReset;
  assign mem_sparse_2_metaReset = metaReset;
  assign io_dataInstr_0_data = {_T_69,_T_68}; // @[memory.scala 82:16]
  assign mem_sparse_clock = clock;
  assign mem_sparse_io_w_1_addr = io_dw_addr;
  assign mem_sparse_io_w_1_en = io_dw_en;
  assign mem_sparse_io_w_1_data = io_dw_data[7:0];
  assign mem_sparse_io_r_0_addr = underlying_0__T_54_addr_pipe_0;
  assign mem_sparse_0_clock = clock;
  assign mem_sparse_0_io_w_1_addr = io_dw_addr;
  assign mem_sparse_0_io_w_1_en = io_dw_en;
  assign mem_sparse_0_io_w_1_data = io_dw_data[15:8];
  assign mem_sparse_0_io_r_0_addr = underlying_1__T_54_addr_pipe_0;
  assign mem_sparse_1_clock = clock;
  assign mem_sparse_1_io_w_1_addr = io_dw_addr;
  assign mem_sparse_1_io_w_1_en = io_dw_en;
  assign mem_sparse_1_io_w_1_data = io_dw_data[23:16];
  assign mem_sparse_1_io_r_0_addr = underlying_2__T_54_addr_pipe_0;
  assign mem_sparse_2_clock = clock;
  assign mem_sparse_2_io_w_1_addr = io_dw_addr;
  assign mem_sparse_2_io_w_1_en = io_dw_en;
  assign mem_sparse_2_io_w_1_data = io_dw_data[31:24];
  assign mem_sparse_2_io_r_0_addr = underlying_3__T_54_addr_pipe_0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  underlying_0__T_54_addr_pipe_0 = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  underlying_1__T_54_addr_pipe_0 = _RAND_1[20:0];
  _RAND_2 = {1{`RANDOM}};
  underlying_2__T_54_addr_pipe_0 = _RAND_2[20:0];
  _RAND_3 = {1{`RANDOM}};
  underlying_3__T_54_addr_pipe_0 = _RAND_3[20:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      underlying_0__T_54_addr_pipe_0 <= 21'h0;
    end else begin
      underlying_0__T_54_addr_pipe_0 <= io_dataInstr_0_addr;
    end
    if (metaReset) begin
      underlying_1__T_54_addr_pipe_0 <= 21'h0;
    end else begin
      underlying_1__T_54_addr_pipe_0 <= io_dataInstr_0_addr;
    end
    if (metaReset) begin
      underlying_2__T_54_addr_pipe_0 <= 21'h0;
    end else begin
      underlying_2__T_54_addr_pipe_0 <= io_dataInstr_0_addr;
    end
    if (metaReset) begin
      underlying_3__T_54_addr_pipe_0 <= 21'h0;
    end else begin
      underlying_3__T_54_addr_pipe_0 <= io_dataInstr_0_addr;
    end
  end
endmodule
module SparseMem_0(
  input         metaReset,
  input         clock,
  input  [20:0] io_w_1_addr,
  input         io_w_1_en,
  input  [7:0]  io_w_1_data,
  input  [20:0] io_r_0_addr,
  output [7:0]  io_r_0_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] mem [0:31];
  wire [7:0] mem__T_152_data;
  wire [4:0] mem__T_152_addr;
  wire [7:0] mem__T_274_data;
  wire [4:0] mem__T_274_addr;
  wire [7:0] mem__T_396_data;
  wire [4:0] mem__T_396_addr;
  wire [7:0] mem__T_528_data;
  wire [4:0] mem__T_528_addr;
  wire  mem__T_528_mask;
  wire  mem__T_528_en;
  wire [7:0] mem__T_656_data;
  wire [4:0] mem__T_656_addr;
  wire  mem__T_656_mask;
  wire  mem__T_656_en;
  reg [20:0] addresses_0_bits;
  reg [20:0] addresses_1_bits;
  reg [20:0] addresses_2_bits;
  reg [20:0] addresses_3_bits;
  reg [20:0] addresses_4_bits;
  reg [20:0] addresses_5_bits;
  reg [20:0] addresses_6_bits;
  reg [20:0] addresses_7_bits;
  reg [20:0] addresses_8_bits;
  reg [20:0] addresses_9_bits;
  reg [20:0] addresses_10_bits;
  reg [20:0] addresses_11_bits;
  reg [20:0] addresses_12_bits;
  reg [20:0] addresses_13_bits;
  reg [20:0] addresses_14_bits;
  reg [20:0] addresses_15_bits;
  reg [20:0] addresses_16_bits;
  reg [20:0] addresses_17_bits;
  reg [20:0] addresses_18_bits;
  reg [20:0] addresses_19_bits;
  reg [20:0] addresses_20_bits;
  reg [20:0] addresses_21_bits;
  reg [20:0] addresses_22_bits;
  reg [20:0] addresses_23_bits;
  reg [20:0] addresses_24_bits;
  reg [20:0] addresses_25_bits;
  reg [20:0] addresses_26_bits;
  reg [20:0] addresses_27_bits;
  reg [20:0] addresses_28_bits;
  reg [20:0] addresses_29_bits;
  reg [20:0] addresses_30_bits;
  reg [20:0] addresses_31_bits;
  wire  _T_33 = addresses_0_bits == io_r_0_addr;
  wire  _T_35 = addresses_1_bits == io_r_0_addr;
  wire  _T_37 = addresses_2_bits == io_r_0_addr;
  wire  _T_39 = addresses_3_bits == io_r_0_addr;
  wire  _T_41 = addresses_4_bits == io_r_0_addr;
  wire  _T_43 = addresses_5_bits == io_r_0_addr;
  wire  _T_45 = addresses_6_bits == io_r_0_addr;
  wire  _T_47 = addresses_7_bits == io_r_0_addr;
  wire  _T_49 = addresses_8_bits == io_r_0_addr;
  wire  _T_51 = addresses_9_bits == io_r_0_addr;
  wire  _T_53 = addresses_10_bits == io_r_0_addr;
  wire  _T_55 = addresses_11_bits == io_r_0_addr;
  wire  _T_57 = addresses_12_bits == io_r_0_addr;
  wire  _T_59 = addresses_13_bits == io_r_0_addr;
  wire  _T_61 = addresses_14_bits == io_r_0_addr;
  wire  _T_63 = addresses_15_bits == io_r_0_addr;
  wire  _T_65 = addresses_16_bits == io_r_0_addr;
  wire  _T_67 = addresses_17_bits == io_r_0_addr;
  wire  _T_69 = addresses_18_bits == io_r_0_addr;
  wire  _T_71 = addresses_19_bits == io_r_0_addr;
  wire  _T_73 = addresses_20_bits == io_r_0_addr;
  wire  _T_75 = addresses_21_bits == io_r_0_addr;
  wire  _T_77 = addresses_22_bits == io_r_0_addr;
  wire  _T_79 = addresses_23_bits == io_r_0_addr;
  wire  _T_81 = addresses_24_bits == io_r_0_addr;
  wire  _T_83 = addresses_25_bits == io_r_0_addr;
  wire  _T_85 = addresses_26_bits == io_r_0_addr;
  wire  _T_87 = addresses_27_bits == io_r_0_addr;
  wire  _T_89 = addresses_28_bits == io_r_0_addr;
  wire  _T_91 = addresses_29_bits == io_r_0_addr;
  wire  _T_93 = addresses_30_bits == io_r_0_addr;
  wire  _T_95 = addresses_31_bits == io_r_0_addr;
  wire [7:0] _T_104 = {_T_47,_T_45,_T_43,_T_41,_T_39,_T_37,_T_35,_T_33};
  wire [15:0] _T_112 = {_T_63,_T_61,_T_59,_T_57,_T_55,_T_53,_T_51,_T_49,_T_104};
  wire [7:0] _T_119 = {_T_79,_T_77,_T_75,_T_73,_T_71,_T_69,_T_67,_T_65};
  wire [31:0] _T_128 = {_T_95,_T_93,_T_91,_T_89,_T_87,_T_85,_T_83,_T_81,_T_119,_T_112};
  wire  _T_129 = _T_128 != 32'h0;
  wire  _T_132 = |_T_128[31:16];
  wire [15:0] _T_133 = _T_128[31:16] | _T_128[15:0];
  wire  _T_136 = |_T_133[15:8];
  wire [7:0] _T_137 = _T_133[15:8] | _T_133[7:0];
  wire  _T_140 = |_T_137[7:4];
  wire [3:0] _T_141 = _T_137[7:4] | _T_137[3:0];
  wire  _T_144 = |_T_141[3:2];
  wire [1:0] _T_145 = _T_141[3:2] | _T_141[1:0];
  wire [3:0] _T_149 = {_T_136,_T_140,_T_144,_T_145[1]};
  wire  _T_155 = addresses_0_bits == 21'h0;
  wire  _T_157 = addresses_1_bits == 21'h0;
  wire  _T_159 = addresses_2_bits == 21'h0;
  wire  _T_161 = addresses_3_bits == 21'h0;
  wire  _T_163 = addresses_4_bits == 21'h0;
  wire  _T_165 = addresses_5_bits == 21'h0;
  wire  _T_167 = addresses_6_bits == 21'h0;
  wire  _T_169 = addresses_7_bits == 21'h0;
  wire  _T_171 = addresses_8_bits == 21'h0;
  wire  _T_173 = addresses_9_bits == 21'h0;
  wire  _T_175 = addresses_10_bits == 21'h0;
  wire  _T_177 = addresses_11_bits == 21'h0;
  wire  _T_179 = addresses_12_bits == 21'h0;
  wire  _T_181 = addresses_13_bits == 21'h0;
  wire  _T_183 = addresses_14_bits == 21'h0;
  wire  _T_185 = addresses_15_bits == 21'h0;
  wire  _T_187 = addresses_16_bits == 21'h0;
  wire  _T_189 = addresses_17_bits == 21'h0;
  wire  _T_191 = addresses_18_bits == 21'h0;
  wire  _T_193 = addresses_19_bits == 21'h0;
  wire  _T_195 = addresses_20_bits == 21'h0;
  wire  _T_197 = addresses_21_bits == 21'h0;
  wire  _T_199 = addresses_22_bits == 21'h0;
  wire  _T_201 = addresses_23_bits == 21'h0;
  wire  _T_203 = addresses_24_bits == 21'h0;
  wire  _T_205 = addresses_25_bits == 21'h0;
  wire  _T_207 = addresses_26_bits == 21'h0;
  wire  _T_209 = addresses_27_bits == 21'h0;
  wire  _T_211 = addresses_28_bits == 21'h0;
  wire  _T_213 = addresses_29_bits == 21'h0;
  wire  _T_215 = addresses_30_bits == 21'h0;
  wire  _T_217 = addresses_31_bits == 21'h0;
  wire [7:0] _T_226 = {_T_169,_T_167,_T_165,_T_163,_T_161,_T_159,_T_157,_T_155};
  wire [15:0] _T_234 = {_T_185,_T_183,_T_181,_T_179,_T_177,_T_175,_T_173,_T_171,_T_226};
  wire [7:0] _T_241 = {_T_201,_T_199,_T_197,_T_195,_T_193,_T_191,_T_189,_T_187};
  wire [31:0] _T_250 = {_T_217,_T_215,_T_213,_T_211,_T_209,_T_207,_T_205,_T_203,_T_241,_T_234};
  wire  _T_251 = _T_250 != 32'h0;
  wire  _T_254 = |_T_250[31:16];
  wire [15:0] _T_255 = _T_250[31:16] | _T_250[15:0];
  wire  _T_258 = |_T_255[15:8];
  wire [7:0] _T_259 = _T_255[15:8] | _T_255[7:0];
  wire  _T_262 = |_T_259[7:4];
  wire [3:0] _T_263 = _T_259[7:4] | _T_259[3:0];
  wire  _T_266 = |_T_263[3:2];
  wire [1:0] _T_267 = _T_263[3:2] | _T_263[1:0];
  wire [3:0] _T_271 = {_T_258,_T_262,_T_266,_T_267[1]};
  wire [4:0] _T_272 = {_T_254,_T_258,_T_262,_T_266,_T_267[1]};
  reg [5:0] nextAddr;
  wire [5:0] _T_400 = nextAddr + 6'h1;
  wire [5:0] _T_524 = _T_251 ? {{1'd0}, _T_272} : nextAddr;
  wire  _T_532 = addresses_0_bits == io_w_1_addr;
  wire  _T_534 = addresses_1_bits == io_w_1_addr;
  wire  _T_536 = addresses_2_bits == io_w_1_addr;
  wire  _T_538 = addresses_3_bits == io_w_1_addr;
  wire  _T_540 = addresses_4_bits == io_w_1_addr;
  wire  _T_542 = addresses_5_bits == io_w_1_addr;
  wire  _T_544 = addresses_6_bits == io_w_1_addr;
  wire  _T_546 = addresses_7_bits == io_w_1_addr;
  wire  _T_548 = addresses_8_bits == io_w_1_addr;
  wire  _T_550 = addresses_9_bits == io_w_1_addr;
  wire  _T_552 = addresses_10_bits == io_w_1_addr;
  wire  _T_554 = addresses_11_bits == io_w_1_addr;
  wire  _T_556 = addresses_12_bits == io_w_1_addr;
  wire  _T_558 = addresses_13_bits == io_w_1_addr;
  wire  _T_560 = addresses_14_bits == io_w_1_addr;
  wire  _T_562 = addresses_15_bits == io_w_1_addr;
  wire  _T_564 = addresses_16_bits == io_w_1_addr;
  wire  _T_566 = addresses_17_bits == io_w_1_addr;
  wire  _T_568 = addresses_18_bits == io_w_1_addr;
  wire  _T_570 = addresses_19_bits == io_w_1_addr;
  wire  _T_572 = addresses_20_bits == io_w_1_addr;
  wire  _T_574 = addresses_21_bits == io_w_1_addr;
  wire  _T_576 = addresses_22_bits == io_w_1_addr;
  wire  _T_578 = addresses_23_bits == io_w_1_addr;
  wire  _T_580 = addresses_24_bits == io_w_1_addr;
  wire  _T_582 = addresses_25_bits == io_w_1_addr;
  wire  _T_584 = addresses_26_bits == io_w_1_addr;
  wire  _T_586 = addresses_27_bits == io_w_1_addr;
  wire  _T_588 = addresses_28_bits == io_w_1_addr;
  wire  _T_590 = addresses_29_bits == io_w_1_addr;
  wire  _T_592 = addresses_30_bits == io_w_1_addr;
  wire  _T_594 = addresses_31_bits == io_w_1_addr;
  wire [7:0] _T_603 = {_T_546,_T_544,_T_542,_T_540,_T_538,_T_536,_T_534,_T_532};
  wire [15:0] _T_611 = {_T_562,_T_560,_T_558,_T_556,_T_554,_T_552,_T_550,_T_548,_T_603};
  wire [7:0] _T_618 = {_T_578,_T_576,_T_574,_T_572,_T_570,_T_568,_T_566,_T_564};
  wire [31:0] _T_627 = {_T_594,_T_592,_T_590,_T_588,_T_586,_T_584,_T_582,_T_580,_T_618,_T_611};
  wire  _T_628 = _T_627 != 32'h0;
  wire  _T_631 = |_T_627[31:16];
  wire [15:0] _T_632 = _T_627[31:16] | _T_627[15:0];
  wire  _T_635 = |_T_632[15:8];
  wire [7:0] _T_636 = _T_632[15:8] | _T_632[7:0];
  wire  _T_639 = |_T_636[7:4];
  wire [3:0] _T_640 = _T_636[7:4] | _T_636[3:0];
  wire  _T_643 = |_T_640[3:2];
  wire [1:0] _T_644 = _T_640[3:2] | _T_640[1:0];
  wire [4:0] _T_649 = {_T_631,_T_635,_T_639,_T_643,_T_644[1]};
  wire  _T_650 = ~_T_628;
  wire  _T_651 = io_w_1_en & _T_650;
  wire [5:0] _T_652 = _T_628 ? {{1'd0}, _T_649} : nextAddr;
  wire [5:0] nextAddrUpdate = _T_651 ? _T_400 : nextAddr;
  wire  _T_659 = nextAddrUpdate <= 6'h20;
  wire  _T_662 = ~_T_659;
  assign mem__T_152_addr = {_T_132,_T_149};
  assign mem__T_152_data = mem[mem__T_152_addr];
  assign mem__T_274_addr = {_T_254,_T_271};
  assign mem__T_274_data = mem[mem__T_274_addr];
  assign mem__T_396_addr = {_T_254,_T_271};
  assign mem__T_396_data = mem[mem__T_396_addr];
  assign mem__T_528_data = 8'h0;
  assign mem__T_528_addr = _T_524[4:0];
  assign mem__T_528_mask = 1'h1;
  assign mem__T_528_en = 1'h0;
  assign mem__T_656_data = io_w_1_data;
  assign mem__T_656_addr = _T_652[4:0];
  assign mem__T_656_mask = 1'h1;
  assign mem__T_656_en = io_w_1_en;
  assign io_r_0_data = _T_129 ? mem__T_152_data : 8'h0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  addresses_0_bits = _RAND_1[20:0];
  _RAND_2 = {1{`RANDOM}};
  addresses_1_bits = _RAND_2[20:0];
  _RAND_3 = {1{`RANDOM}};
  addresses_2_bits = _RAND_3[20:0];
  _RAND_4 = {1{`RANDOM}};
  addresses_3_bits = _RAND_4[20:0];
  _RAND_5 = {1{`RANDOM}};
  addresses_4_bits = _RAND_5[20:0];
  _RAND_6 = {1{`RANDOM}};
  addresses_5_bits = _RAND_6[20:0];
  _RAND_7 = {1{`RANDOM}};
  addresses_6_bits = _RAND_7[20:0];
  _RAND_8 = {1{`RANDOM}};
  addresses_7_bits = _RAND_8[20:0];
  _RAND_9 = {1{`RANDOM}};
  addresses_8_bits = _RAND_9[20:0];
  _RAND_10 = {1{`RANDOM}};
  addresses_9_bits = _RAND_10[20:0];
  _RAND_11 = {1{`RANDOM}};
  addresses_10_bits = _RAND_11[20:0];
  _RAND_12 = {1{`RANDOM}};
  addresses_11_bits = _RAND_12[20:0];
  _RAND_13 = {1{`RANDOM}};
  addresses_12_bits = _RAND_13[20:0];
  _RAND_14 = {1{`RANDOM}};
  addresses_13_bits = _RAND_14[20:0];
  _RAND_15 = {1{`RANDOM}};
  addresses_14_bits = _RAND_15[20:0];
  _RAND_16 = {1{`RANDOM}};
  addresses_15_bits = _RAND_16[20:0];
  _RAND_17 = {1{`RANDOM}};
  addresses_16_bits = _RAND_17[20:0];
  _RAND_18 = {1{`RANDOM}};
  addresses_17_bits = _RAND_18[20:0];
  _RAND_19 = {1{`RANDOM}};
  addresses_18_bits = _RAND_19[20:0];
  _RAND_20 = {1{`RANDOM}};
  addresses_19_bits = _RAND_20[20:0];
  _RAND_21 = {1{`RANDOM}};
  addresses_20_bits = _RAND_21[20:0];
  _RAND_22 = {1{`RANDOM}};
  addresses_21_bits = _RAND_22[20:0];
  _RAND_23 = {1{`RANDOM}};
  addresses_22_bits = _RAND_23[20:0];
  _RAND_24 = {1{`RANDOM}};
  addresses_23_bits = _RAND_24[20:0];
  _RAND_25 = {1{`RANDOM}};
  addresses_24_bits = _RAND_25[20:0];
  _RAND_26 = {1{`RANDOM}};
  addresses_25_bits = _RAND_26[20:0];
  _RAND_27 = {1{`RANDOM}};
  addresses_26_bits = _RAND_27[20:0];
  _RAND_28 = {1{`RANDOM}};
  addresses_27_bits = _RAND_28[20:0];
  _RAND_29 = {1{`RANDOM}};
  addresses_28_bits = _RAND_29[20:0];
  _RAND_30 = {1{`RANDOM}};
  addresses_29_bits = _RAND_30[20:0];
  _RAND_31 = {1{`RANDOM}};
  addresses_30_bits = _RAND_31[20:0];
  _RAND_32 = {1{`RANDOM}};
  addresses_31_bits = _RAND_32[20:0];
  _RAND_33 = {1{`RANDOM}};
  nextAddr = _RAND_33[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_528_en & mem__T_528_mask) begin
      mem[mem__T_528_addr] <= mem__T_528_data;
    end
    if(mem__T_656_en & mem__T_656_mask) begin
      mem[mem__T_656_addr] <= mem__T_656_data;
    end
    if (metaReset) begin
      addresses_0_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h0 == _T_652[4:0]) begin
        addresses_0_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_1_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h1 == _T_652[4:0]) begin
        addresses_1_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_2_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h2 == _T_652[4:0]) begin
        addresses_2_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_3_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h3 == _T_652[4:0]) begin
        addresses_3_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_4_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h4 == _T_652[4:0]) begin
        addresses_4_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_5_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h5 == _T_652[4:0]) begin
        addresses_5_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_6_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h6 == _T_652[4:0]) begin
        addresses_6_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_7_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h7 == _T_652[4:0]) begin
        addresses_7_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_8_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h8 == _T_652[4:0]) begin
        addresses_8_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_9_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h9 == _T_652[4:0]) begin
        addresses_9_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_10_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'ha == _T_652[4:0]) begin
        addresses_10_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_11_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'hb == _T_652[4:0]) begin
        addresses_11_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_12_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'hc == _T_652[4:0]) begin
        addresses_12_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_13_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'hd == _T_652[4:0]) begin
        addresses_13_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_14_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'he == _T_652[4:0]) begin
        addresses_14_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_15_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'hf == _T_652[4:0]) begin
        addresses_15_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_16_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h10 == _T_652[4:0]) begin
        addresses_16_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_17_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h11 == _T_652[4:0]) begin
        addresses_17_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_18_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h12 == _T_652[4:0]) begin
        addresses_18_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_19_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h13 == _T_652[4:0]) begin
        addresses_19_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_20_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h14 == _T_652[4:0]) begin
        addresses_20_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_21_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h15 == _T_652[4:0]) begin
        addresses_21_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_22_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h16 == _T_652[4:0]) begin
        addresses_22_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_23_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h17 == _T_652[4:0]) begin
        addresses_23_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_24_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h18 == _T_652[4:0]) begin
        addresses_24_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_25_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h19 == _T_652[4:0]) begin
        addresses_25_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_26_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h1a == _T_652[4:0]) begin
        addresses_26_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_27_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h1b == _T_652[4:0]) begin
        addresses_27_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_28_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h1c == _T_652[4:0]) begin
        addresses_28_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_29_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h1d == _T_652[4:0]) begin
        addresses_29_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_30_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h1e == _T_652[4:0]) begin
        addresses_30_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      addresses_31_bits <= 21'h0;
    end else if (io_w_1_en) begin
      if (5'h1f == _T_652[4:0]) begin
        addresses_31_bits <= io_w_1_addr;
      end
    end
    if (metaReset) begin
      nextAddr <= 6'h0;
    end else if (_T_651) begin
      nextAddr <= _T_400;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_662) begin
          $fwrite(32'h80000002,"Assertion failed: SparseMem ran out of space with size %d, increase size in ReplaceMemsTransform!\n    at SparseMem.scala:102 assert(nextAddrUpdate <= depth.U,\n",6'h20);
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_662) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SyncScratchPadMemory(
  input         metaReset,
  input         clock,
  input  [31:0] io_core_ports_0_req_bits_addr,
  input  [31:0] io_core_ports_0_req_bits_data,
  input         io_core_ports_0_req_bits_fcn,
  input  [2:0]  io_core_ports_0_req_bits_typ,
  output [31:0] io_core_ports_0_resp_bits_data,
  output        _GEN_1_0,
  output        _GEN_4_0,
  output        _GEN_0_1,
  output        _GEN_3_1,
  output        _GEN_2_1,
  output        _GEN_5_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  sync_data_metaReset; // @[memory.scala 199:26]
  wire  sync_data_clock; // @[memory.scala 199:26]
  wire [20:0] sync_data_io_dataInstr_0_addr; // @[memory.scala 199:26]
  wire [31:0] sync_data_io_dataInstr_0_data; // @[memory.scala 199:26]
  wire [20:0] sync_data_io_dw_addr; // @[memory.scala 199:26]
  wire [31:0] sync_data_io_dw_data; // @[memory.scala 199:26]
  wire  sync_data_io_dw_en; // @[memory.scala 199:26]
  reg [2:0] req_typi; // @[memory.scala 213:22]
  wire  _T_233 = req_typi == 3'h1; // @[memory.scala 218:17]
  wire [23:0] _T_238 = sync_data_io_dataInstr_0_data[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_240 = {_T_238,sync_data_io_dataInstr_0_data[7:0]}; // @[Cat.scala 30:58]
  wire  _T_241 = req_typi == 3'h2; // @[memory.scala 219:17]
  wire [15:0] _T_246 = sync_data_io_dataInstr_0_data[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_248 = {_T_246,sync_data_io_dataInstr_0_data[15:0]}; // @[Cat.scala 30:58]
  wire  _T_249 = req_typi == 3'h5; // @[memory.scala 220:17]
  wire [31:0] _T_256 = {24'h0,sync_data_io_dataInstr_0_data[7:0]}; // @[Cat.scala 30:58]
  wire  _T_257 = req_typi == 3'h6; // @[memory.scala 221:17]
  wire [31:0] _T_264 = {16'h0,sync_data_io_dataInstr_0_data[15:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_265 = _T_257 ? _T_264 : sync_data_io_dataInstr_0_data; // @[Mux.scala 61:16]
  wire [31:0] _T_266 = _T_249 ? _T_256 : _T_265; // @[Mux.scala 61:16]
  wire [31:0] _T_267 = _T_241 ? _T_248 : _T_266; // @[Mux.scala 61:16]
  wire [4:0] _T_276 = {io_core_ports_0_req_bits_addr[1:0], 3'h0}; // @[memory.scala 227:85]
  wire [62:0] _GEN_8 = {{31'd0}, io_core_ports_0_req_bits_data}; // @[memory.scala 227:66]
  wire [62:0] _T_277 = _GEN_8 << _T_276; // @[memory.scala 227:66]
  wire [31:0] _T_280 = {io_core_ports_0_req_bits_addr[31:2],2'h0}; // @[Cat.scala 30:58]
  SyncMem sync_data ( // @[memory.scala 199:26]
    .metaReset(sync_data_metaReset),
    .clock(sync_data_clock),
    .io_dataInstr_0_addr(sync_data_io_dataInstr_0_addr),
    .io_dataInstr_0_data(sync_data_io_dataInstr_0_data),
    .io_dw_addr(sync_data_io_dw_addr),
    .io_dw_data(sync_data_io_dw_data),
    .io_dw_en(sync_data_io_dw_en)
  );
  assign sync_data_metaReset = metaReset;
  assign io_core_ports_0_resp_bits_data = _T_233 ? _T_240 : _T_267; // @[memory.scala 217:40]
  assign _GEN_1_0 = sync_data_io_dataInstr_0_data[15];
  assign _GEN_4_0 = req_typi == 3'h2;
  assign _GEN_0_1 = sync_data_io_dataInstr_0_data[7];
  assign _GEN_3_1 = req_typi == 3'h5;
  assign _GEN_2_1 = req_typi == 3'h6;
  assign _GEN_5_1 = req_typi == 3'h1;
  assign sync_data_clock = clock;
  assign sync_data_io_dataInstr_0_addr = io_core_ports_0_req_bits_addr[20:0]; // @[memory.scala 206:38]
  assign sync_data_io_dw_addr = _T_280[20:0]; // @[memory.scala 228:28]
  assign sync_data_io_dw_data = _T_277[31:0]; // @[memory.scala 227:28]
  assign sync_data_io_dw_en = io_core_ports_0_req_bits_fcn; // @[memory.scala 224:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  req_typi = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (metaReset) begin
      req_typi <= 3'h0;
    end else begin
      req_typi <= io_core_ports_0_req_bits_typ;
    end
  end
endmodule
